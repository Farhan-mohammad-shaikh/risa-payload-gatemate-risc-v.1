//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 January 2025)
//  Compile Time: 1970-01-01 00:59:59
//  Program Run:  2025-02-27 00:39:15
//  Program Call: p_r +uCIO -ccf colognechip_gatemate_evb.ccf -cCP -A 1 -i colognechip_gatemate_evb_synth.v -o colognechip_gatemate_evb -lib ccag 
//  File Type:    Verilog

// Gatecount:   7303
module colognechip_gatemate_evb (cdone_ice40 , clk10 , power_fauld_ice40 , spi_flash_miso , spi_ice40_miso , uart_ice40_rx , 
       uart_logging_rx , usb_uart_rx ,
       core_en_ice40 , hyperram_clk_n , hyperram_clk_p , hyperram_cs_n , hyperram_rst_n , osc_en_ice40 , 
       spi_flash_clk , spi_flash_cs_n , spi_flash_mosi , spi_ice40_clk , spi_ice40_cs_n , spi_ice40_mosi , 
       uart_ice40_tx , uart_logging_tx , usb_uart_tx , user_led_n0 , user_led_n1 , user_led_n2 , 
       user_led_n3 , vio_en_ice40 ,
       creset_ice40 , gatemate_debug_3 , gatemate_debug_4 , gatemate_debug_5 , hyperram_dq , hyperram_rwds , 
       i2c0_scl , i2c0_sda , i2c1_scl , i2c1_sda , ice40_io_vcore_0 , ice40_io_vcore_1 , 
       ice40_io_vcore_2 , ice40_io_vcore_4 , ice40_io_vio_0 , ice40_io_vio_1 , ice40_io_vio_2 , ice40_io_vio_3 , 
       ice40_io_vio_4 , ice40_io_vio_5 
) ;

input  cdone_ice40;
input  clk10;
input  power_fauld_ice40;
input  spi_flash_miso;
input  spi_ice40_miso;
input  uart_ice40_rx;
input  uart_logging_rx;
input  usb_uart_rx;

output core_en_ice40;
output hyperram_clk_n;
output hyperram_clk_p;
output hyperram_cs_n;
output hyperram_rst_n;
output osc_en_ice40;
output spi_flash_clk;
output spi_flash_cs_n;
output spi_flash_mosi;
output spi_ice40_clk;
output spi_ice40_cs_n;
output spi_ice40_mosi;
output uart_ice40_tx;
output uart_logging_tx;
output usb_uart_tx;
output user_led_n0;
output user_led_n1;
output user_led_n2;
output user_led_n3;
output vio_en_ice40;

inout  creset_ice40;
inout  gatemate_debug_3;
inout  gatemate_debug_4;
inout  gatemate_debug_5;
inout  [7:0]hyperram_dq;
inout  hyperram_rwds;
inout  i2c0_scl;
inout  i2c0_sda;
inout  i2c1_scl;
inout  i2c1_sda;
inout  ice40_io_vcore_0;
inout  ice40_io_vcore_1;
inout  ice40_io_vcore_2;
inout  ice40_io_vcore_4;
inout  ice40_io_vio_0;
inout  ice40_io_vio_1;
inout  ice40_io_vio_2;
inout  ice40_io_vio_3;
inout  ice40_io_vio_4;
inout  ice40_io_vio_5;


wire [7:0]hyperram_dq;
wire clk10;
wire na1_1;
wire na2_1;
wire na3_1;
wire na4_2;
wire na5_1;
wire na6_2;
wire na8_1;
wire na8_2;
wire na9_1;
wire na12_1;
wire na13_1;
wire na15_1;
wire na16_1;
wire na17_1;
wire na18_1;
wire na19_1;
wire na20_1;
wire na21_1;
wire na22_1;
wire na23_1;
wire na24_1;
wire na25_1;
wire na26_2;
wire na27_1;
wire na28_1;
wire na29_1;
wire na30_1;
wire na31_2;
wire na32_1;
wire na34_2;
wire na35_1;
wire na36_1;
wire na36_2;
wire na37_1;
wire na39_1;
wire na41_1;
wire na42_2;
wire na43_1;
wire na43_2;
wire na45_1;
wire na46_1;
wire na46_1_i;
wire na47_2;
wire na48_1;
wire na50_1;
wire na50_2;
wire na51_1;
wire na53_1;
wire na55_1;
wire na56_2;
wire na57_1;
wire na58_1;
wire na58_1_i;
wire na59_1;
wire na61_1;
wire na63_1;
wire na64_1;
wire na66_1;
wire na67_1;
wire na67_2;
wire na68_2;
wire na69_1;
wire na70_1;
wire na71_1;
wire na72_1;
wire na73_1;
wire na74_1;
wire na75_1;
wire na76_2;
wire na77_2;
wire na78_1;
wire na79_1;
wire na80_1;
wire na81_1;
wire na81_2;
wire na82_1;
wire na83_1;
wire na83_1_i;
wire na84_1;
wire na85_1;
wire na86_1;
wire na87_1;
wire na88_1;
wire na88_2;
wire na89_1;
wire na89_2;
wire na90_1;
wire na90_2;
wire na91_1;
wire na91_2;
wire na92_1;
wire na92_2;
wire na95_1;
wire na95_2;
wire na97_1;
wire na97_2;
wire na99_2;
wire na100_2;
wire na101_2;
wire na102_1;
wire na103_1;
wire na103_2;
wire na104_1;
wire na106_1;
wire na106_2;
wire na107_1;
wire na107_2;
wire na112_2;
wire na114_1;
wire na116_1;
wire na116_2;
wire na120_2;
wire na122_1;
wire na125_1;
wire na128_1;
wire na129_1;
wire na129_2;
wire na133_1;
wire na135_1;
wire na135_2;
wire na138_1;
wire na140_1;
wire na142_1;
wire na142_2;
wire na144_1;
wire na145_1;
wire na147_1;
wire na149_1;
wire na149_2;
wire na151_1;
wire na152_1;
wire na154_1;
wire na154_2;
wire na155_1;
wire na157_1;
wire na159_1;
wire na159_2;
wire na160_1;
wire na160_1_i;
wire na161_2;
wire na164_1;
wire na164_1_i;
wire na165_1;
wire na165_1_i;
wire na166_1;
wire na166_1_i;
wire na167_1;
wire na167_1_i;
wire na168_1;
wire na168_1_i;
wire na169_2;
wire na170_1;
wire na170_1_i;
wire na171_1;
wire na171_1_i;
wire na172_2;
wire na173_1;
wire na174_1;
wire na177_1;
wire na178_2;
wire na179_1;
wire na180_1;
wire na180_2;
wire na182_1;
wire na186_1;
wire na189_1;
wire na193_1;
wire na194_1;
wire na197_1;
wire na199_1;
wire na203_1;
wire na207_1;
wire na210_1;
wire na211_2;
wire na212_1;
wire na214_1;
wire na214_2;
wire na215_1;
wire na220_1;
wire na223_1;
wire na224_1;
wire na228_1;
wire na232_1;
wire na232_2;
wire na233_1;
wire na234_2;
wire na235_1;
wire na235_1_i;
wire na236_1;
wire na236_2;
wire na237_1;
wire na238_2;
wire na239_1;
wire na239_2;
wire na240_1;
wire na240_2;
wire na241_1;
wire na241_2;
wire na242_1;
wire na242_2;
wire na243_1;
wire na243_2;
wire na244_1;
wire na244_2;
wire na245_1;
wire na245_2;
wire na246_1;
wire na246_1_i;
wire na247_1;
wire na247_1_i;
wire na248_2;
wire na251_1;
wire na251_2;
wire na252_1;
wire na254_1;
wire na256_2;
wire na257_1;
wire na258_2;
wire na259_1;
wire na259_2;
wire na260_1;
wire na260_2;
wire na261_1;
wire na261_2;
wire na262_1;
wire na262_2;
wire na263_1;
wire na263_2;
wire na264_1;
wire na264_2;
wire na265_1;
wire na265_2;
wire na266_1;
wire na266_1_i;
wire na267_1;
wire na267_1_i;
wire na268_1;
wire na269_1;
wire na269_1_i;
wire na270_1;
wire na270_1_i;
wire na271_1;
wire na271_1_i;
wire na272_1;
wire na272_1_i;
wire na273_1;
wire na277_1;
wire na278_1;
wire na279_1;
wire na279_1_i;
wire na280_2;
wire na281_2;
wire na281_2_i;
wire na282_1;
wire na282_1_i;
wire na283_2;
wire na285_1;
wire na287_1;
wire na288_2;
wire na289_1;
wire na289_1_i;
wire na289_2;
wire na289_2_i;
wire na290_1;
wire na291_1;
wire na291_1_i;
wire na291_2;
wire na291_2_i;
wire na292_1;
wire na294_1;
wire na295_1;
wire na295_1_i;
wire na296_1;
wire na298_1;
wire na298_2;
wire na299_2;
wire na300_1;
wire na300_1_i;
wire na301_2;
wire na301_2_i;
wire na303_1;
wire na306_1;
wire na306_1_i;
wire na307_2;
wire na308_1;
wire na309_1;
wire na309_1_i;
wire na310_1;
wire na311_1;
wire na311_1_i;
wire na312_2;
wire na313_1;
wire na313_1_i;
wire na316_1;
wire na318_1;
wire na318_1_i;
wire na318_2;
wire na318_2_i;
wire na320_1;
wire na320_1_i;
wire na320_2;
wire na320_2_i;
wire na321_2;
wire na321_2_i;
wire na322_1;
wire na322_1_i;
wire na324_1;
wire na325_1;
wire na325_2;
wire na326_2;
wire na326_2_i;
wire na329_1;
wire na331_1;
wire na332_2;
wire na333_1;
wire na333_1_i;
wire na334_1;
wire na334_1_i;
wire na335_1;
wire na336_1;
wire na336_1_i;
wire na336_2;
wire na336_2_i;
wire na337_1;
wire na338_2;
wire na338_2_i;
wire na339_1;
wire na340_1;
wire na341_1;
wire na343_1;
wire na344_2;
wire na346_1;
wire na346_2;
wire na347_1;
wire na347_2;
wire na348_1;
wire na349_1;
wire na350_1;
wire na351_1;
wire na353_1;
wire na353_2;
wire na354_1;
wire na354_2;
wire na355_1;
wire na356_1;
wire na356_2;
wire na357_1;
wire na358_1;
wire na359_1;
wire na359_2;
wire na364_2;
wire na365_2;
wire na369_1;
wire na369_2;
wire na374_1;
wire na378_1;
wire na378_2;
wire na379_1;
wire na380_2;
wire na383_2;
wire na385_1;
wire na386_1;
wire na387_2;
wire na389_1;
wire na389_2;
wire na393_2;
wire na396_1;
wire na397_2;
wire na399_1;
wire na401_2;
wire na401_2_i;
wire na402_1;
wire na403_1;
wire na403_2;
wire na404_1;
wire na404_1_i;
wire na404_2;
wire na404_2_i;
wire na406_1;
wire na406_2;
wire na407_2;
wire na408_1;
wire na408_1_i;
wire na409_1;
wire na410_1;
wire na412_2;
wire na412_2_i;
wire na413_1;
wire na413_1_i;
wire na414_2;
wire na414_2_i;
wire na415_1;
wire na415_1_i;
wire na416_1;
wire na416_1_i;
wire na417_1;
wire na417_1_i;
wire na418_1;
wire na418_1_i;
wire na419_1;
wire na419_1_i;
wire na420_1;
wire na420_1_i;
wire na421_1;
wire na423_1;
wire na423_1_i;
wire na424_1;
wire na424_1_i;
wire na425_1;
wire na425_1_i;
wire na426_2;
wire na427_2;
wire na428_1;
wire na428_2;
wire na429_2;
wire na430_1;
wire na431_1;
wire na432_1;
wire na433_1;
wire na433_2;
wire na435_1;
wire na435_2;
wire na436_1;
wire na437_1;
wire na437_1_i;
wire na438_1;
wire na438_1_i;
wire na439_1;
wire na439_1_i;
wire na440_1;
wire na440_1_i;
wire na441_1;
wire na441_1_i;
wire na442_1;
wire na442_1_i;
wire na443_1;
wire na443_1_i;
wire na444_1;
wire na445_1;
wire na445_1_i;
wire na446_1;
wire na446_1_i;
wire na447_1;
wire na447_1_i;
wire na448_1;
wire na450_2;
wire na452_1;
wire na452_2;
wire na454_1;
wire na454_2;
wire na455_1;
wire na455_1_i;
wire na456_1;
wire na456_1_i;
wire na457_1;
wire na457_1_i;
wire na459_1;
wire na463_1;
wire na463_2;
wire na464_1;
wire na464_1_i;
wire na467_1;
wire na468_1;
wire na469_1;
wire na469_2;
wire na470_1;
wire na470_1_i;
wire na471_1;
wire na471_1_i;
wire na472_1;
wire na473_1;
wire na473_1_i;
wire na474_1;
wire na474_1_i;
wire na475_1;
wire na475_1_i;
wire na476_1;
wire na476_1_i;
wire na477_1;
wire na477_1_i;
wire na478_1;
wire na478_2;
wire na479_1;
wire na479_1_i;
wire na480_1;
wire na480_1_i;
wire na481_1;
wire na481_1_i;
wire na482_2;
wire na483_1;
wire na483_1_i;
wire na484_1;
wire na484_1_i;
wire na485_1;
wire na485_1_i;
wire na486_1;
wire na486_1_i;
wire na488_1;
wire na488_2;
wire na489_1;
wire na490_2;
wire na492_1;
wire na492_1_i;
wire na493_1;
wire na493_1_i;
wire na494_1;
wire na494_1_i;
wire na495_1;
wire na495_1_i;
wire na496_1;
wire na496_1_i;
wire na497_1;
wire na497_1_i;
wire na498_1;
wire na498_1_i;
wire na498_2;
wire na498_2_i;
wire na499_2;
wire na500_1;
wire na500_2;
wire na501_1;
wire na501_1_i;
wire na502_2;
wire na503_2;
wire na504_1;
wire na505_1;
wire na505_1_i;
wire na505_2;
wire na505_2_i;
wire na506_2;
wire na507_1;
wire na507_1_i;
wire na508_1;
wire na511_1;
wire na511_2;
wire na514_2;
wire na515_1;
wire na515_1_i;
wire na516_1;
wire na517_1;
wire na517_1_i;
wire na517_2;
wire na517_2_i;
wire na520_1;
wire na520_2;
wire na521_1;
wire na521_1_i;
wire na522_2;
wire na523_1;
wire na523_1_i;
wire na526_2;
wire na527_1;
wire na528_1;
wire na531_1;
wire na531_1_i;
wire na531_2;
wire na531_2_i;
wire na532_1;
wire na533_1;
wire na536_1;
wire na536_2;
wire na537_1;
wire na540_1;
wire na542_1;
wire na542_2;
wire na545_1;
wire na546_1;
wire na546_1_i;
wire na546_2;
wire na546_2_i;
wire na547_1;
wire na547_2;
wire na548_1;
wire na550_1;
wire na551_1;
wire na551_1_i;
wire na552_1;
wire na552_2;
wire na554_2;
wire na555_1;
wire na557_2;
wire na557_2_i;
wire na558_1;
wire na558_1_i;
wire na560_1;
wire na560_1_i;
wire na561_1;
wire na561_1_i;
wire na561_2;
wire na561_2_i;
wire na562_2;
wire na563_1;
wire na563_1_i;
wire na564_1;
wire na565_2;
wire na566_1;
wire na567_1;
wire na568_1;
wire na568_1_i;
wire na569_2;
wire na570_1;
wire na570_1_i;
wire na571_1;
wire na571_1_i;
wire na572_1;
wire na573_1;
wire na573_1_i;
wire na574_1;
wire na574_2;
wire na576_1;
wire na578_1;
wire na578_1_i;
wire na579_1;
wire na579_1_i;
wire na581_1;
wire na581_2;
wire na582_1;
wire na582_2;
wire na584_1;
wire na587_1;
wire na587_1_i;
wire na587_2;
wire na587_2_i;
wire na588_1;
wire na588_2;
wire na589_1;
wire na589_2;
wire na590_1;
wire na592_2;
wire na592_2_i;
wire na593_1;
wire na593_2;
wire na594_1;
wire na595_1;
wire na597_1;
wire na597_1_i;
wire na598_1;
wire na598_2;
wire na600_1;
wire na602_2;
wire na602_2_i;
wire na603_1;
wire na603_2;
wire na604_1;
wire na607_1;
wire na608_1;
wire na608_1_i;
wire na609_1;
wire na609_2;
wire na610_1;
wire na612_1;
wire na613_2;
wire na613_2_i;
wire na614_1;
wire na614_2;
wire na615_1;
wire na617_1;
wire na618_1;
wire na618_1_i;
wire na619_1;
wire na619_2;
wire na620_1;
wire na622_1;
wire na623_2;
wire na623_2_i;
wire na624_1;
wire na624_2;
wire na625_1;
wire na627_1;
wire na628_1;
wire na628_1_i;
wire na629_1;
wire na629_2;
wire na630_1;
wire na632_1;
wire na633_2;
wire na633_2_i;
wire na634_1;
wire na634_2;
wire na635_1;
wire na637_1;
wire na638_1;
wire na638_1_i;
wire na639_1;
wire na639_1_i;
wire na640_2;
wire na640_2_i;
wire na641_1;
wire na641_1_i;
wire na643_1;
wire na647_1;
wire na649_2;
wire na650_1;
wire na652_1;
wire na652_2;
wire na654_1;
wire na655_1;
wire na656_1;
wire na657_1;
wire na658_1;
wire na658_2;
wire na659_1;
wire na661_1;
wire na662_2;
wire na662_2_i;
wire na663_1;
wire na663_1_i;
wire na664_1;
wire na664_2;
wire na665_1;
wire na667_1;
wire na668_1;
wire na668_1_i;
wire na669_1;
wire na669_2;
wire na670_1;
wire na672_1;
wire na673_2;
wire na673_2_i;
wire na674_1;
wire na674_2;
wire na675_1;
wire na677_1;
wire na678_1;
wire na678_1_i;
wire na679_1;
wire na679_2;
wire na680_1;
wire na682_1;
wire na683_2;
wire na683_2_i;
wire na684_1;
wire na684_2;
wire na685_1;
wire na687_1;
wire na688_1;
wire na688_1_i;
wire na689_1;
wire na689_2;
wire na690_1;
wire na692_1;
wire na693_2;
wire na693_2_i;
wire na694_1;
wire na694_2;
wire na695_1;
wire na697_1;
wire na698_1;
wire na698_1_i;
wire na699_1;
wire na699_2;
wire na700_1;
wire na702_1;
wire na703_2;
wire na703_2_i;
wire na704_1;
wire na704_2;
wire na705_1;
wire na707_1;
wire na708_2;
wire na708_2_i;
wire na709_1;
wire na709_1_i;
wire na709_2;
wire na709_2_i;
wire na710_1;
wire na711_1;
wire na712_1;
wire na712_1_i;
wire na713_1;
wire na714_1;
wire na714_2;
wire na716_1;
wire na718_1;
wire na718_2;
wire na719_1;
wire na719_2;
wire na720_1;
wire na723_1;
wire na724_1;
wire na724_1_i;
wire na725_1;
wire na725_1_i;
wire na727_2;
wire na728_1;
wire na728_2;
wire na729_1;
wire na730_1;
wire na731_1;
wire na734_2;
wire na736_2;
wire na737_1;
wire na737_2;
wire na738_1;
wire na739_1;
wire na740_1;
wire na740_1_i;
wire na740_2;
wire na740_2_i;
wire na741_1;
wire na741_2;
wire na742_1;
wire na743_1;
wire na745_1;
wire na745_2;
wire na746_1;
wire na747_1;
wire na748_1;
wire na748_1_i;
wire na748_2;
wire na748_2_i;
wire na749_1;
wire na749_2;
wire na750_1;
wire na751_1;
wire na753_1;
wire na753_1_i;
wire na753_2;
wire na753_2_i;
wire na754_1;
wire na755_2;
wire na755_2_i;
wire na756_1;
wire na757_1;
wire na757_1_i;
wire na758_1;
wire na758_2;
wire na759_1;
wire na759_2;
wire na760_1;
wire na761_1;
wire na763_1;
wire na763_2;
wire na764_1;
wire na765_1;
wire na766_1;
wire na766_1_i;
wire na766_2;
wire na766_2_i;
wire na767_1;
wire na767_2;
wire na768_1;
wire na769_1;
wire na771_1;
wire na771_2;
wire na772_1;
wire na773_1;
wire na774_1;
wire na774_1_i;
wire na774_2;
wire na774_2_i;
wire na775_1;
wire na775_2;
wire na776_1;
wire na777_1;
wire na779_1;
wire na779_2;
wire na780_1;
wire na781_1;
wire na782_1;
wire na782_1_i;
wire na782_2;
wire na782_2_i;
wire na783_1;
wire na783_1_i;
wire na784_2;
wire na785_1;
wire na785_1_i;
wire na786_1;
wire na786_2;
wire na787_1;
wire na788_1;
wire na790_2;
wire na790_2_i;
wire na791_1;
wire na791_1_i;
wire na792_1;
wire na792_2;
wire na793_1;
wire na794_1;
wire na795_1;
wire na795_1_i;
wire na795_2;
wire na795_2_i;
wire na796_1;
wire na796_1_i;
wire na797_1;
wire na798_2;
wire na799_1;
wire na799_2;
wire na800_1;
wire na801_1;
wire na803_1;
wire na803_2;
wire na804_1;
wire na805_1;
wire na806_1;
wire na806_1_i;
wire na806_2;
wire na806_2_i;
wire na807_1;
wire na807_2;
wire na808_1;
wire na809_1;
wire na810_1;
wire na810_1_i;
wire na810_2;
wire na810_2_i;
wire na811_1;
wire na811_2;
wire na812_1;
wire na813_1;
wire na815_1;
wire na815_2;
wire na816_1;
wire na817_1;
wire na819_1;
wire na819_2;
wire na820_1;
wire na821_1;
wire na822_1;
wire na822_1_i;
wire na822_2;
wire na822_2_i;
wire na823_1;
wire na823_2;
wire na824_1;
wire na825_1;
wire na826_1;
wire na826_1_i;
wire na826_2;
wire na826_2_i;
wire na827_1;
wire na827_1_i;
wire na828_1;
wire na828_2;
wire na829_1;
wire na830_1;
wire na831_1;
wire na831_1_i;
wire na831_2;
wire na831_2_i;
wire na832_1;
wire na832_1_i;
wire na833_1;
wire na834_1;
wire na834_2;
wire na835_1;
wire na836_1;
wire na838_1;
wire na838_1_i;
wire na839_1;
wire na839_1_i;
wire na841_2;
wire na843_1;
wire na843_2;
wire na844_1;
wire na845_1;
wire na847_1;
wire na847_2;
wire na848_1;
wire na849_1;
wire na851_2;
wire na851_2_i;
wire na853_2;
wire na854_1;
wire na855_1;
wire na856_2;
wire na857_1;
wire na857_2;
wire na858_1;
wire na859_1;
wire na860_1;
wire na860_1_i;
wire na860_2;
wire na860_2_i;
wire na861_2;
wire na861_2_i;
wire na863_1;
wire na863_2;
wire na864_1;
wire na865_1;
wire na866_1;
wire na866_1_i;
wire na866_2;
wire na866_2_i;
wire na867_1;
wire na867_1_i;
wire na868_1;
wire na868_1_i;
wire na869_1;
wire na869_1_i;
wire na870_1;
wire na870_1_i;
wire na870_2;
wire na870_2_i;
wire na871_2;
wire na872_1;
wire na872_1_i;
wire na873_2;
wire na874_1;
wire na875_1;
wire na875_1_i;
wire na876_1;
wire na877_1;
wire na877_1_i;
wire na878_1;
wire na878_1_i;
wire na878_2;
wire na878_2_i;
wire na879_1;
wire na879_1_i;
wire na880_1;
wire na880_1_i;
wire na881_1;
wire na881_1_i;
wire na882_1;
wire na882_1_i;
wire na883_1;
wire na883_1_i;
wire na884_1;
wire na884_1_i;
wire na886_1;
wire na886_1_i;
wire na888_2;
wire na888_2_i;
wire na890_1;
wire na890_1_i;
wire na891_1;
wire na891_1_i;
wire na892_1;
wire na892_1_i;
wire na893_2;
wire na894_1;
wire na894_1_i;
wire na895_1;
wire na895_1_i;
wire na896_1;
wire na896_1_i;
wire na897_1;
wire na897_1_i;
wire na898_1;
wire na900_1;
wire na900_1_i;
wire na901_1;
wire na902_1;
wire na902_1_i;
wire na903_1;
wire na903_1_i;
wire na904_1;
wire na904_1_i;
wire na905_1;
wire na906_1;
wire na907_2;
wire na907_2_i;
wire na908_1;
wire na909_1;
wire na909_1_i;
wire na911_2;
wire na911_2_i;
wire na912_1;
wire na912_1_i;
wire na913_1;
wire na913_1_i;
wire na913_2;
wire na913_2_i;
wire na914_1;
wire na915_2;
wire na916_1;
wire na916_1_i;
wire na917_1;
wire na917_1_i;
wire na918_1;
wire na918_1_i;
wire na919_1;
wire na919_1_i;
wire na920_1;
wire na920_1_i;
wire na921_1;
wire na921_1_i;
wire na923_1;
wire na924_1;
wire na925_1;
wire na925_1_i;
wire na925_2;
wire na925_2_i;
wire na926_1;
wire na927_2;
wire na927_2_i;
wire na928_1;
wire na929_2;
wire na930_1;
wire na930_1_i;
wire na931_1;
wire na932_1;
wire na933_1;
wire na933_1_i;
wire na934_2;
wire na935_1;
wire na935_1_i;
wire na936_1;
wire na936_1_i;
wire na937_1;
wire na937_1_i;
wire na938_1;
wire na938_1_i;
wire na939_1;
wire na939_1_i;
wire na940_1;
wire na940_1_i;
wire na941_1;
wire na941_1_i;
wire na942_1;
wire na942_1_i;
wire na943_1;
wire na944_1;
wire na945_1;
wire na945_1_i;
wire na946_2;
wire na947_1;
wire na948_1;
wire na948_1_i;
wire na949_1;
wire na949_1_i;
wire na950_1;
wire na950_1_i;
wire na950_2;
wire na950_2_i;
wire na951_1;
wire na951_2;
wire na952_1;
wire na952_1_i;
wire na952_2;
wire na952_2_i;
wire na953_1;
wire na953_1_i;
wire na954_1;
wire na955_1;
wire na957_1;
wire na957_1_i;
wire na957_2;
wire na957_2_i;
wire na958_1;
wire na958_1_i;
wire na959_1;
wire na959_1_i;
wire na959_2;
wire na959_2_i;
wire na960_1;
wire na960_1_i;
wire na961_2;
wire na962_1;
wire na962_1_i;
wire na963_1;
wire na963_1_i;
wire na964_1;
wire na964_1_i;
wire na964_2;
wire na964_2_i;
wire na965_1;
wire na965_1_i;
wire na965_2;
wire na965_2_i;
wire na966_1;
wire na966_1_i;
wire na966_2;
wire na966_2_i;
wire na967_1;
wire na967_1_i;
wire na967_2;
wire na967_2_i;
wire na968_1;
wire na968_1_i;
wire na968_2;
wire na968_2_i;
wire na969_1;
wire na969_1_i;
wire na969_2;
wire na969_2_i;
wire na970_1;
wire na970_1_i;
wire na970_2;
wire na970_2_i;
wire na971_1;
wire na971_1_i;
wire na973_1;
wire na973_1_i;
wire na974_1;
wire na977_1;
wire na977_1_i;
wire na977_2;
wire na977_2_i;
wire na978_1;
wire na978_1_i;
wire na979_1;
wire na979_1_i;
wire na980_1;
wire na980_1_i;
wire na981_1;
wire na981_1_i;
wire na983_1;
wire na984_1;
wire na984_1_i;
wire na984_2;
wire na984_2_i;
wire na985_1;
wire na985_1_i;
wire na985_2;
wire na985_2_i;
wire na986_1;
wire na988_1;
wire na989_1;
wire na990_1;
wire na990_1_i;
wire na991_2;
wire na992_1;
wire na992_1_i;
wire na993_1;
wire na995_1;
wire na995_1_i;
wire na996_2;
wire na997_1;
wire na998_1;
wire na999_1;
wire na999_1_i;
wire na999_2;
wire na999_2_i;
wire i2c0_scl;
wire i2c0_sda;
wire i2c1_scl;
wire i2c1_sda;
wire na1000_1;
wire na1000_1_i;
wire na1001_1;
wire na1001_1_i;
wire na1002_1;
wire na1002_1_i;
wire na1003_1;
wire na1003_1_i;
wire na1004_1;
wire na1004_1_i;
wire na1005_1;
wire na1005_1_i;
wire na1006_2;
wire na1006_2_i;
wire na1007_1;
wire na1007_1_i;
wire na1008_2;
wire na1008_2_i;
wire na1009_1;
wire na1009_1_i;
wire na1010_1;
wire na1010_1_i;
wire na1011_2;
wire na1012_1;
wire na1013_1;
wire na1013_2;
wire na1014_2;
wire na1016_1;
wire na1016_1_i;
wire na1017_1;
wire na1018_1;
wire na1018_1_i;
wire na1019_1;
wire na1020_1;
wire na1020_1_i;
wire na1021_1;
wire na1021_1_i;
wire na1022_1;
wire na1022_1_i;
wire na1023_1;
wire na1024_1;
wire na1026_1;
wire na1026_1_i;
wire na1027_1;
wire na1028_1;
wire na1030_1;
wire na1030_1_i;
wire na1032_1;
wire na1032_1_i;
wire na1033_1;
wire na1033_1_i;
wire na1034_1;
wire na1034_2;
wire na1035_1;
wire na1035_1_i;
wire na1036_2;
wire na1036_2_i;
wire na1037_2;
wire na1038_1;
wire na1038_1_i;
wire na1038_2;
wire na1038_2_i;
wire na1039_1;
wire na1039_1_i;
wire na1040_1;
wire na1040_1_i;
wire na1042_1;
wire na1045_2;
wire na1046_2;
wire na1048_2;
wire na1048_2_i;
wire na1049_1;
wire na1053_1;
wire na1053_1_i;
wire na1053_2;
wire na1053_2_i;
wire na1054_2;
wire na1055_1;
wire na1057_1;
wire na1057_1_i;
wire na1057_2;
wire na1057_2_i;
wire na1059_1;
wire na1059_1_i;
wire na1059_2;
wire na1059_2_i;
wire na1061_1;
wire na1061_1_i;
wire na1061_2;
wire na1061_2_i;
wire na1062_1;
wire na1063_1;
wire na1064_1;
wire na1064_1_i;
wire na1064_2;
wire na1064_2_i;
wire na1065_1;
wire na1065_1_i;
wire na1065_2;
wire na1065_2_i;
wire na1066_1;
wire na1067_2;
wire na1068_1;
wire na1068_1_i;
wire na1069_1;
wire na1069_1_i;
wire na1070_1;
wire na1070_1_i;
wire na1071_1;
wire na1071_1_i;
wire na1072_1;
wire na1072_1_i;
wire na1073_1;
wire na1073_2;
wire na1074_1;
wire na1074_1_i;
wire na1075_1;
wire na1075_1_i;
wire na1076_1;
wire na1076_1_i;
wire na1077_1;
wire na1077_1_i;
wire na1078_1;
wire na1079_1;
wire na1079_1_i;
wire na1080_1;
wire na1080_1_i;
wire na1081_1;
wire na1081_1_i;
wire na1082_1;
wire na1082_1_i;
wire na1083_1;
wire na1083_1_i;
wire na1084_1;
wire na1084_1_i;
wire na1085_1;
wire na1085_1_i;
wire na1086_1;
wire na1086_1_i;
wire na1087_1;
wire na1087_1_i;
wire na1088_1;
wire na1088_1_i;
wire na1089_1;
wire na1089_1_i;
wire na1090_1;
wire na1090_1_i;
wire na1091_1;
wire na1092_1;
wire na1092_1_i;
wire na1093_1;
wire na1093_1_i;
wire na1094_1;
wire na1094_1_i;
wire na1095_2;
wire na1096_1;
wire na1096_1_i;
wire na1097_2;
wire na1098_1;
wire na1098_1_i;
wire na1099_1;
wire na1100_1;
wire na1100_1_i;
wire na1101_2;
wire na1102_1;
wire na1102_1_i;
wire na1103_1;
wire na1104_1;
wire na1104_1_i;
wire na1105_2;
wire na1106_1;
wire na1106_1_i;
wire na1108_1;
wire na1109_1;
wire na1109_1_i;
wire na1110_1;
wire na1111_1;
wire na1111_1_i;
wire na1112_2;
wire na1113_1;
wire na1113_1_i;
wire na1113_2;
wire na1113_2_i;
wire na1114_1;
wire na1114_1_i;
wire na1115_1;
wire na1115_1_i;
wire na1116_1;
wire na1116_1_i;
wire na1117_1;
wire na1117_1_i;
wire na1118_1;
wire na1118_1_i;
wire na1119_1;
wire na1119_1_i;
wire na1120_1;
wire na1121_1;
wire na1121_1_i;
wire na1123_1;
wire na1123_1_i;
wire na1124_1;
wire na1124_1_i;
wire na1125_2;
wire na1125_2_i;
wire na1126_1;
wire na1126_1_i;
wire na1126_2;
wire na1126_2_i;
wire na1127_1;
wire na1127_1_i;
wire na1128_2;
wire na1128_2_i;
wire na1129_1;
wire na1130_1;
wire na1130_2;
wire na1131_1;
wire na1132_1;
wire na1134_1;
wire na1134_1_i;
wire na1134_2;
wire na1134_2_i;
wire na1135_1;
wire na1136_2;
wire na1137_1;
wire na1138_1;
wire na1138_1_i;
wire na1139_1;
wire na1140_1;
wire na1140_1_i;
wire na1141_1;
wire na1142_1;
wire na1142_1_i;
wire na1143_2;
wire na1145_1;
wire na1145_1_i;
wire na1147_1;
wire na1147_1_i;
wire na1148_1;
wire na1148_1_i;
wire na1149_1;
wire na1149_1_i;
wire na1150_1;
wire na1150_1_i;
wire na1151_1;
wire na1151_1_i;
wire na1152_1;
wire na1152_1_i;
wire na1153_1;
wire na1153_1_i;
wire na1154_1;
wire na1154_1_i;
wire na1155_1;
wire na1155_1_i;
wire na1156_1;
wire na1156_1_i;
wire na1157_1;
wire na1157_1_i;
wire na1158_1;
wire na1158_1_i;
wire na1159_1;
wire na1159_1_i;
wire na1160_1;
wire na1160_2;
wire na1161_1;
wire na1161_1_i;
wire na1162_1;
wire na1162_1_i;
wire na1163_1;
wire na1163_1_i;
wire na1164_1;
wire na1164_1_i;
wire na1165_1;
wire na1165_1_i;
wire na1165_2;
wire na1165_2_i;
wire na1166_1;
wire na1167_1;
wire na1167_1_i;
wire na1168_1;
wire na1169_1;
wire na1169_1_i;
wire na1170_1;
wire na1170_1_i;
wire na1171_1;
wire na1171_1_i;
wire na1172_1;
wire na1172_1_i;
wire na1173_1;
wire na1173_1_i;
wire na1174_2;
wire na1175_1;
wire na1175_1_i;
wire na1175_2;
wire na1175_2_i;
wire na1176_2;
wire na1177_1;
wire na1177_1_i;
wire na1177_2;
wire na1177_2_i;
wire na1178_2;
wire na1179_1;
wire na1181_1;
wire na1181_2;
wire na1182_1;
wire na1184_1;
wire na1184_1_i;
wire na1185_1;
wire na1185_1_i;
wire na1186_1;
wire na1186_1_i;
wire na1187_1;
wire na1187_1_i;
wire na1188_1;
wire na1188_1_i;
wire na1189_2;
wire na1190_1;
wire na1191_1;
wire na1191_1_i;
wire na1191_2;
wire na1191_2_i;
wire na1192_1;
wire na1193_1;
wire na1193_1_i;
wire na1193_2;
wire na1193_2_i;
wire na1194_1;
wire na1196_1;
wire na1197_1;
wire na1197_1_i;
wire na1198_1;
wire na1198_1_i;
wire na1199_1;
wire na1199_1_i;
wire na1200_1;
wire na1200_1_i;
wire na1201_1;
wire na1201_1_i;
wire na1202_1;
wire na1202_1_i;
wire na1203_1;
wire na1203_1_i;
wire na1204_1;
wire na1204_1_i;
wire na1205_1;
wire na1205_1_i;
wire na1206_1;
wire na1206_1_i;
wire na1207_1;
wire na1207_1_i;
wire na1208_1;
wire na1208_1_i;
wire na1209_1;
wire na1209_1_i;
wire na1210_1;
wire na1210_1_i;
wire na1211_1;
wire na1212_2;
wire na1212_2_i;
wire na1213_1;
wire na1213_1_i;
wire na1214_1;
wire na1215_1;
wire na1215_1_i;
wire na1216_1;
wire na1216_1_i;
wire na1218_2;
wire na1219_1;
wire na1219_1_i;
wire na1220_1;
wire na1220_1_i;
wire na1221_1;
wire na1221_1_i;
wire na1222_1;
wire na1222_1_i;
wire na1223_1;
wire na1223_1_i;
wire na1224_1;
wire na1224_1_i;
wire na1225_1;
wire na1225_1_i;
wire na1226_1;
wire na1226_1_i;
wire na1227_1;
wire na1227_1_i;
wire na1228_1;
wire na1228_1_i;
wire na1229_1;
wire na1229_1_i;
wire na1230_1;
wire na1230_1_i;
wire na1231_1;
wire na1231_1_i;
wire na1232_1;
wire na1232_1_i;
wire na1233_1;
wire na1233_1_i;
wire na1234_1;
wire na1234_1_i;
wire na1236_1;
wire na1237_1;
wire na1238_1;
wire na1238_1_i;
wire na1239_1;
wire na1239_1_i;
wire na1240_1;
wire na1240_1_i;
wire na1241_1;
wire na1241_1_i;
wire na1242_1;
wire na1242_1_i;
wire na1243_1;
wire na1243_1_i;
wire na1244_1;
wire na1244_1_i;
wire na1245_1;
wire na1245_1_i;
wire na1246_1;
wire na1246_1_i;
wire na1247_2;
wire na1248_1;
wire na1248_1_i;
wire na1249_1;
wire na1249_1_i;
wire na1250_1;
wire na1250_1_i;
wire na1250_2;
wire na1250_2_i;
wire na1252_1;
wire na1252_1_i;
wire na1252_2;
wire na1252_2_i;
wire na1254_1;
wire na1254_1_i;
wire na1254_2;
wire na1254_2_i;
wire na1256_1;
wire na1256_1_i;
wire na1256_2;
wire na1256_2_i;
wire na1258_1;
wire na1258_1_i;
wire na1258_2;
wire na1258_2_i;
wire na1260_1;
wire na1260_1_i;
wire na1260_2;
wire na1260_2_i;
wire na1261_1;
wire na1261_1_i;
wire na1262_1;
wire na1262_1_i;
wire na1263_1;
wire na1263_1_i;
wire na1264_1;
wire na1264_1_i;
wire na1265_1;
wire na1265_1_i;
wire na1266_1;
wire na1266_1_i;
wire na1267_1;
wire na1267_1_i;
wire na1268_1;
wire na1268_1_i;
wire na1269_1;
wire na1269_1_i;
wire na1270_1;
wire na1270_1_i;
wire na1271_1;
wire na1271_1_i;
wire na1272_1;
wire na1272_1_i;
wire na1273_1;
wire na1273_1_i;
wire na1274_1;
wire na1274_1_i;
wire na1275_1;
wire na1279_1;
wire na1281_2;
wire na1282_1;
wire na1283_2;
wire na1284_1;
wire na1284_2;
wire na1285_1;
wire na1286_2;
wire na1287_1;
wire na1287_1_i;
wire na1288_1;
wire na1289_1;
wire na1289_1_i;
wire na1290_1;
wire na1291_1;
wire na1291_1_i;
wire na1292_1;
wire na1293_1;
wire na1293_1_i;
wire na1294_1;
wire na1295_1;
wire na1295_1_i;
wire na1296_1;
wire na1297_1;
wire na1297_1_i;
wire na1298_1;
wire na1299_1;
wire na1299_1_i;
wire na1300_1;
wire na1301_1;
wire na1301_1_i;
wire na1302_1;
wire na1303_1;
wire na1303_1_i;
wire na1304_1;
wire na1306_1;
wire na1307_2;
wire na1308_1;
wire na1308_1_i;
wire na1309_1;
wire na1310_1;
wire na1310_1_i;
wire na1311_1;
wire na1312_1;
wire na1312_1_i;
wire na1313_1;
wire na1314_1;
wire na1314_1_i;
wire na1314_2;
wire na1314_2_i;
wire na1315_1;
wire na1316_1;
wire na1316_1_i;
wire na1317_1;
wire na1318_1;
wire na1318_1_i;
wire na1319_1;
wire na1321_1;
wire na1322_1;
wire na1323_1;
wire na1323_1_i;
wire na1324_1;
wire na1325_1;
wire na1325_1_i;
wire na1326_1;
wire na1327_1;
wire na1327_1_i;
wire na1328_1;
wire na1329_1;
wire na1329_1_i;
wire na1330_1;
wire na1331_1;
wire na1331_1_i;
wire na1332_1;
wire na1333_1;
wire na1333_1_i;
wire na1334_1;
wire na1335_1;
wire na1335_1_i;
wire na1336_1;
wire na1337_1;
wire na1337_1_i;
wire na1337_2;
wire na1337_2_i;
wire na1338_1;
wire na1339_1;
wire na1340_1;
wire na1340_1_i;
wire na1341_1;
wire na1342_1;
wire na1342_1_i;
wire na1343_1;
wire na1343_1_i;
wire na1343_2;
wire na1343_2_i;
wire na1344_2;
wire na1344_2_i;
wire na1345_1;
wire na1346_1;
wire na1346_1_i;
wire na1347_1;
wire na1349_2;
wire na1349_2_i;
wire na1350_1;
wire na1350_1_i;
wire na1351_1;
wire na1351_1_i;
wire na1352_1;
wire na1353_1;
wire na1353_1_i;
wire na1354_1;
wire na1354_1_i;
wire na1355_1;
wire na1355_1_i;
wire na1355_2;
wire na1355_2_i;
wire na1356_1;
wire na1357_2;
wire na1358_1;
wire na1358_1_i;
wire na1359_1;
wire na1359_1_i;
wire na1359_2;
wire na1359_2_i;
wire na1360_1;
wire na1361_1;
wire na1362_1;
wire na1362_1_i;
wire na1363_1;
wire na1363_1_i;
wire na1364_1;
wire na1364_1_i;
wire na1365_1;
wire na1365_1_i;
wire na1365_2;
wire na1365_2_i;
wire na1366_1;
wire na1366_1_i;
wire na1367_1;
wire na1367_1_i;
wire na1370_1;
wire na1370_2;
wire na1371_1;
wire na1371_1_i;
wire na1372_1;
wire na1372_1_i;
wire na1373_2;
wire na1373_2_i;
wire na1375_1;
wire na1375_1_i;
wire na1375_2;
wire na1375_2_i;
wire na1377_1;
wire na1377_1_i;
wire na1378_1;
wire na1379_2;
wire na1379_2_i;
wire na1380_1;
wire na1381_1;
wire na1382_1;
wire na1382_1_i;
wire na1383_1;
wire na1383_1_i;
wire na1384_1;
wire na1385_2;
wire na1387_1;
wire na1387_1_i;
wire na1387_2;
wire na1387_2_i;
wire na1388_1;
wire na1388_1_i;
wire na1389_1;
wire na1390_2;
wire na1390_2_i;
wire na1392_1;
wire na1392_1_i;
wire na1393_1;
wire na1393_2;
wire na1395_1;
wire na1399_2;
wire na1399_2_i;
wire na1400_1;
wire na1401_2;
wire na1401_2_i;
wire na1403_1;
wire na1403_1_i;
wire na1405_1;
wire na1405_1_i;
wire na1407_1;
wire na1407_1_i;
wire na1408_1;
wire na1408_1_i;
wire na1409_1;
wire na1409_1_i;
wire na1411_1;
wire na1411_1_i;
wire na1412_2;
wire na1412_2_i;
wire na1414_2;
wire na1414_2_i;
wire na1415_1;
wire na1415_1_i;
wire na1416_2;
wire na1418_1;
wire na1418_1_i;
wire na1419_1;
wire na1419_1_i;
wire na1420_2;
wire na1420_2_i;
wire na1421_1;
wire na1425_2;
wire na1427_1;
wire na1427_1_i;
wire na1427_2;
wire na1427_2_i;
wire na1429_1;
wire na1429_1_i;
wire na1429_2;
wire na1429_2_i;
wire na1430_1;
wire na1430_1_i;
wire na1431_2;
wire na1431_2_i;
wire na1433_1;
wire na1433_1_i;
wire na1433_2;
wire na1433_2_i;
wire na1434_2;
wire na1435_1;
wire na1435_1_i;
wire na1436_1;
wire na1438_1;
wire na1438_1_i;
wire na1441_1;
wire na1441_1_i;
wire na1443_2;
wire na1443_2_i;
wire na1445_1;
wire na1445_1_i;
wire na1446_1;
wire na1447_1;
wire na1451_1;
wire na1453_1;
wire na1454_2;
wire na1455_1;
wire na1456_1;
wire na1456_2;
wire na1457_2;
wire na1458_1;
wire na1458_1_i;
wire na1460_2;
wire na1460_2_i;
wire na1462_1;
wire na1462_1_i;
wire na1462_2;
wire na1462_2_i;
wire na1463_2;
wire na1464_2;
wire na1464_2_i;
wire na1467_1;
wire na1470_2;
wire na1470_2_i;
wire na1471_1;
wire na1473_2;
wire na1473_2_i;
wire na1475_1;
wire na1475_1_i;
wire na1476_1;
wire na1479_1;
wire na1479_1_i;
wire na1481_1;
wire na1481_1_i;
wire na1481_2;
wire na1481_2_i;
wire na1482_1;
wire na1482_1_i;
wire na1484_2;
wire na1484_2_i;
wire na1486_1;
wire na1486_1_i;
wire na1488_2;
wire na1488_2_i;
wire na1490_1;
wire na1490_1_i;
wire na1492_1;
wire na1492_1_i;
wire na1493_1;
wire na1494_1;
wire na1494_2;
wire na1495_1;
wire na1496_1;
wire na1497_1;
wire na1497_1_i;
wire na1497_2;
wire na1497_2_i;
wire na1498_1;
wire na1498_2;
wire na1499_1;
wire na1500_1;
wire na1502_1;
wire na1502_2;
wire na1503_1;
wire na1504_1;
wire na1506_2;
wire na1506_2_i;
wire na1509_1;
wire na1509_1_i;
wire na1512_1;
wire na1512_1_i;
wire na1524_1;
wire na1525_1;
wire na1525_2;
wire na1527_1;
wire na1530_1;
wire na1531_1;
wire na1532_1;
wire na1532_1_i;
wire na1535_1;
wire na1535_1_i;
wire na1538_2;
wire na1538_2_i;
wire na1542_1;
wire na1542_1_i;
wire na1545_2;
wire na1545_2_i;
wire na1548_2;
wire na1548_2_i;
wire na1550_2;
wire na1550_2_i;
wire na1552_1;
wire na1552_2;
wire na1553_1;
wire na1554_1;
wire na1555_1;
wire na1555_1_i;
wire na1555_2;
wire na1555_2_i;
wire na1556_2;
wire na1556_2_i;
wire na1558_2;
wire na1558_2_i;
wire na1560_2;
wire na1560_2_i;
wire na1562_2;
wire na1562_2_i;
wire na1564_2;
wire na1564_2_i;
wire na1568_2;
wire na1568_2_i;
wire na1571_2;
wire na1571_2_i;
wire na1573_1;
wire na1573_1_i;
wire na1575_1;
wire na1575_1_i;
wire na1577_2;
wire na1577_2_i;
wire na1579_2;
wire na1579_2_i;
wire na1583_1;
wire na1583_2;
wire na1584_1;
wire na1586_1;
wire na1587_1;
wire na1587_1_i;
wire na1590_2;
wire na1590_2_i;
wire na1595_2;
wire na1597_1;
wire na1597_1_i;
wire na1598_1;
wire na1599_1;
wire na1599_1_i;
wire na1599_2;
wire na1599_2_i;
wire na1600_1;
wire na1600_2;
wire na1601_1;
wire na1603_1;
wire na1604_1;
wire na1604_1_i;
wire na1605_1;
wire na1605_1_i;
wire na1605_2;
wire na1605_2_i;
wire na1606_1;
wire na1606_1_i;
wire na1606_2;
wire na1606_2_i;
wire na1607_1;
wire na1607_1_i;
wire na1607_2;
wire na1607_2_i;
wire na1612_1;
wire na1614_1;
wire na1616_1;
wire na1616_1_i;
wire na1618_2;
wire na1618_2_i;
wire na1620_1;
wire na1620_1_i;
wire na1621_2;
wire na1621_2_i;
wire na1623_1;
wire na1623_1_i;
wire na1624_1;
wire na1624_1_i;
wire na1626_2;
wire na1626_2_i;
wire na1627_1;
wire na1627_1_i;
wire na1629_2;
wire na1629_2_i;
wire na1631_1;
wire na1631_1_i;
wire na1633_2;
wire na1633_2_i;
wire na1635_2;
wire na1635_2_i;
wire na1637_1;
wire na1637_1_i;
wire na1639_1;
wire na1639_1_i;
wire na1641_2;
wire na1641_2_i;
wire na1643_1;
wire na1643_1_i;
wire na1645_2;
wire na1645_2_i;
wire na1647_2;
wire na1647_2_i;
wire na1649_2;
wire na1649_2_i;
wire na1651_1;
wire na1651_1_i;
wire na1653_1;
wire na1653_1_i;
wire na1654_1;
wire na1654_1_i;
wire na1656_1;
wire na1656_1_i;
wire na1658_1;
wire na1658_1_i;
wire na1659_1;
wire na1659_1_i;
wire na1661_2;
wire na1661_2_i;
wire na1663_1;
wire na1663_1_i;
wire na1665_2;
wire na1665_2_i;
wire na1667_1;
wire na1667_1_i;
wire na1669_2;
wire na1669_2_i;
wire na1677_2;
wire na1677_2_i;
wire na1679_1;
wire na1679_1_i;
wire na1679_2;
wire na1679_2_i;
wire na1681_1;
wire na1681_1_i;
wire na1681_2;
wire na1681_2_i;
wire na1683_1;
wire na1683_1_i;
wire na1683_2;
wire na1683_2_i;
wire na1684_1;
wire na1689_2;
wire na1689_2_i;
wire na1691_1;
wire na1691_1_i;
wire na1693_1;
wire na1693_1_i;
wire na1694_1;
wire na1694_1_i;
wire na1695_1;
wire na1695_1_i;
wire na1697_1;
wire na1697_1_i;
wire na1698_2;
wire na1698_2_i;
wire na1700_1;
wire na1700_1_i;
wire na1702_2;
wire na1702_2_i;
wire na1704_2;
wire na1704_2_i;
wire na1706_2;
wire na1706_2_i;
wire na1708_1;
wire na1708_1_i;
wire na1710_2;
wire na1710_2_i;
wire na1712_1;
wire na1712_1_i;
wire na1714_2;
wire na1714_2_i;
wire na1716_2;
wire na1716_2_i;
wire na1718_2;
wire na1718_2_i;
wire na1720_1;
wire na1720_1_i;
wire na1722_2;
wire na1722_2_i;
wire na1724_1;
wire na1724_1_i;
wire na1726_1;
wire na1726_1_i;
wire na1727_1;
wire na1727_1_i;
wire na1728_1;
wire na1729_2;
wire na1730_1;
wire na1731_2;
wire na1731_2_i;
wire na1733_2;
wire na1733_2_i;
wire na1735_1;
wire na1735_1_i;
wire na1737_1;
wire na1737_1_i;
wire na1739_2;
wire na1739_2_i;
wire na1741_1;
wire na1741_1_i;
wire na1743_1;
wire na1743_1_i;
wire na1743_2;
wire na1743_2_i;
wire na1745_1;
wire na1745_1_i;
wire na1745_2;
wire na1745_2_i;
wire na1747_1;
wire na1747_1_i;
wire na1747_2;
wire na1747_2_i;
wire na1749_1;
wire na1749_1_i;
wire na1749_2;
wire na1749_2_i;
wire na1750_1;
wire na1755_2;
wire na1755_2_i;
wire na1758_1;
wire na1758_1_i;
wire na1761_1;
wire na1761_1_i;
wire na1762_2;
wire na1764_2;
wire na1764_2_i;
wire na1766_2;
wire na1766_2_i;
wire na1768_1;
wire na1768_1_i;
wire na1770_1;
wire na1770_1_i;
wire na1770_2;
wire na1770_2_i;
wire na1774_1;
wire na1774_1_i;
wire na1774_2;
wire na1774_2_i;
wire na1776_1;
wire na1776_1_i;
wire na1780_1;
wire na1780_1_i;
wire na1783_1;
wire na1783_1_i;
wire na1786_2;
wire na1786_2_i;
wire na1792_1;
wire na1792_1_i;
wire na1792_2;
wire na1792_2_i;
wire na1795_2;
wire na1795_2_i;
wire na1798_2;
wire na1798_2_i;
wire na1801_2;
wire na1801_2_i;
wire na1803_1;
wire na1803_1_i;
wire na1804_2;
wire na1804_2_i;
wire na1806_2;
wire na1806_2_i;
wire na1808_1;
wire na1808_1_i;
wire na1810_2;
wire na1810_2_i;
wire na1812_2;
wire na1812_2_i;
wire na1814_1;
wire na1814_1_i;
wire na1816_2;
wire na1816_2_i;
wire na1818_1;
wire na1818_1_i;
wire na1820_1;
wire na1820_1_i;
wire na1822_2;
wire na1822_2_i;
wire na1824_2;
wire na1824_2_i;
wire na1826_2;
wire na1826_2_i;
wire na1828_1;
wire na1828_1_i;
wire na1829_1;
wire na1829_1_i;
wire na1830_2;
wire na1830_2_i;
wire na1832_2;
wire na1832_2_i;
wire na1834_1;
wire na1834_1_i;
wire na1836_2;
wire na1836_2_i;
wire na1838_1;
wire na1838_1_i;
wire na1840_1;
wire na1840_1_i;
wire na1840_2;
wire na1840_2_i;
wire na1842_2;
wire na1842_2_i;
wire na1844_1;
wire na1844_1_i;
wire na1846_2;
wire na1846_2_i;
wire na1848_2;
wire na1848_2_i;
wire na1850_1;
wire na1850_1_i;
wire na1852_2;
wire na1852_2_i;
wire na1854_1;
wire na1854_1_i;
wire na1855_1;
wire na1855_1_i;
wire na1856_1;
wire na1856_1_i;
wire na1858_1;
wire na1858_1_i;
wire na1859_1;
wire na1859_1_i;
wire na1859_2;
wire na1859_2_i;
wire na1860_1;
wire na1860_1_i;
wire na1861_2;
wire na1861_2_i;
wire na1863_1;
wire na1863_1_i;
wire na1864_1;
wire na1864_1_i;
wire na1864_2;
wire na1864_2_i;
wire na1865_1;
wire na1866_1;
wire na1867_1;
wire na1867_1_i;
wire na1868_1;
wire na1868_1_i;
wire na1869_1;
wire na1869_1_i;
wire na1870_1;
wire na1870_1_i;
wire na1872_1;
wire na1875_1;
wire na1877_1;
wire na1879_1;
wire na1880_2;
wire na1880_2_i;
wire na1881_1;
wire na1882_1;
wire na1883_1;
wire na1883_1_i;
wire na1885_1;
wire na1885_1_i;
wire na1886_1;
wire na1886_1_i;
wire na1888_1;
wire na1888_1_i;
wire na1888_2;
wire na1888_2_i;
wire na1889_1;
wire na1889_1_i;
wire na1891_1;
wire na1891_1_i;
wire na1892_1;
wire na1892_1_i;
wire na1893_1;
wire na1893_1_i;
wire na1894_1;
wire na1894_1_i;
wire na1895_2;
wire na1895_2_i;
wire na1896_1;
wire na1897_1;
wire na1897_1_i;
wire na1898_1;
wire na1898_1_i;
wire na1899_1;
wire na1899_1_i;
wire na1900_1;
wire na1900_1_i;
wire na1901_1;
wire na1901_1_i;
wire na1902_1;
wire na1903_1;
wire na1903_1_i;
wire na1904_1;
wire na1904_2;
wire na1905_1;
wire na1907_1;
wire na1909_1;
wire na1910_2;
wire na1911_2;
wire na1914_1;
wire na1914_2;
wire na1915_1;
wire na1915_2;
wire na1917_1;
wire na1918_1;
wire na1920_2;
wire na1921_1;
wire na1921_2;
wire na1922_1;
wire na1922_2;
wire na1927_2;
wire na1929_1;
wire na1930_1;
wire na1930_2;
wire na1931_1;
wire na1932_1;
wire na1932_2;
wire na1937_1;
wire na1939_1;
wire na1940_1;
wire na1940_2;
wire na1941_1;
wire na1942_1;
wire na1942_2;
wire na1944_2;
wire na1949_1;
wire na1949_2;
wire na1950_1;
wire na1951_1;
wire na1951_2;
wire na1953_2;
wire na1958_1;
wire na1958_2;
wire na1959_1;
wire na1960_1;
wire na1960_2;
wire na1962_2;
wire na1967_1;
wire na1967_2;
wire na1968_1;
wire na1969_1;
wire na1969_2;
wire na1971_2;
wire na1976_1;
wire na1976_2;
wire na1977_1;
wire na1978_1;
wire na1978_2;
wire na1980_1;
wire na1981_1;
wire na1982_1;
wire na1984_1;
wire na1986_2;
wire na1987_1;
wire na1987_2;
wire na1990_1;
wire na1990_2;
wire na1991_2;
wire na1993_1;
wire na1994_1;
wire na1994_2;
wire na1997_1;
wire na1997_2;
wire na1998_1;
wire na2000_1;
wire na2001_1;
wire na2001_2;
wire na2004_1;
wire na2004_2;
wire na2005_2;
wire na2007_1;
wire na2008_1;
wire na2008_2;
wire na2011_1;
wire na2011_2;
wire na2012_2;
wire na2014_1;
wire na2015_1;
wire na2015_2;
wire na2018_1;
wire na2018_2;
wire na2019_2;
wire na2021_1;
wire na2022_1;
wire na2022_2;
wire na2025_1;
wire na2025_2;
wire na2026_1;
wire na2028_1;
wire na2029_1;
wire na2029_2;
wire na2032_1;
wire na2032_2;
wire na2033_1;
wire na2035_1;
wire na2036_1;
wire na2036_2;
wire na2039_1;
wire na2039_2;
wire na2040_1;
wire na2042_1;
wire na2043_1;
wire na2043_2;
wire na2045_1;
wire na2045_2;
wire na2046_1;
wire na2047_1;
wire na2048_1;
wire na2050_1;
wire na2050_2;
wire na2052_1;
wire na2052_2;
wire na2053_2;
wire na2054_1;
wire na2055_1;
wire na2057_1;
wire na2057_2;
wire na2059_1;
wire na2059_2;
wire na2060_2;
wire na2061_1;
wire na2062_1;
wire na2064_1;
wire na2064_2;
wire na2066_1;
wire na2066_2;
wire na2067_2;
wire na2068_1;
wire na2069_2;
wire na2071_1;
wire na2071_2;
wire na2073_1;
wire na2073_2;
wire na2074_1;
wire na2075_1;
wire na2076_2;
wire na2078_1;
wire na2078_2;
wire na2080_1;
wire na2080_2;
wire na2081_1;
wire na2082_1;
wire na2083_1;
wire na2085_1;
wire na2085_2;
wire na2087_1;
wire na2087_2;
wire na2088_2;
wire na2089_1;
wire na2090_2;
wire na2092_1;
wire na2092_2;
wire na2094_1;
wire na2094_2;
wire na2095_1;
wire na2096_1;
wire na2097_1;
wire na2099_1;
wire na2099_2;
wire na2101_1;
wire na2101_2;
wire na2102_1;
wire na2103_1;
wire na2104_2;
wire na2106_1;
wire na2106_2;
wire na2108_1;
wire na2108_2;
wire na2109_1;
wire na2110_1;
wire na2111_1;
wire na2113_1;
wire na2113_2;
wire na2115_1;
wire na2115_2;
wire na2116_1;
wire na2117_1;
wire na2118_1;
wire na2120_1;
wire na2120_2;
wire na2122_1;
wire na2122_2;
wire na2123_2;
wire na2124_1;
wire na2125_1;
wire na2127_1;
wire na2127_2;
wire na2129_1;
wire na2129_2;
wire na2130_2;
wire na2131_1;
wire na2132_1;
wire na2134_1;
wire na2134_2;
wire na2136_1;
wire na2136_2;
wire na2137_2;
wire na2138_1;
wire na2139_1;
wire na2141_1;
wire na2141_2;
wire na2143_1;
wire na2143_2;
wire na2144_1;
wire na2145_1;
wire na2146_1;
wire na2148_1;
wire na2148_2;
wire na2150_1;
wire na2150_2;
wire na2151_2;
wire na2152_1;
wire na2153_1;
wire na2155_2;
wire na2155_2_i;
wire na2156_1;
wire na2156_1_i;
wire na2157_1;
wire na2157_1_i;
wire na2158_1;
wire na2158_1_i;
wire na2158_2;
wire na2158_2_i;
wire na2159_1;
wire na2159_1_i;
wire na2160_1;
wire na2161_1;
wire na2161_1_i;
wire na2162_1;
wire na2163_1;
wire na2163_1_i;
wire na2164_2;
wire na2165_1;
wire na2165_1_i;
wire na2166_1;
wire na2166_1_i;
wire na2167_1;
wire na2168_1;
wire na2168_1_i;
wire na2170_1;
wire na2170_1_i;
wire na2171_1;
wire na2171_1_i;
wire na2172_1;
wire na2172_2;
wire na2173_1;
wire na2173_1_i;
wire na2174_2;
wire na2175_1;
wire na2175_1_i;
wire na2176_1;
wire na2177_1;
wire na2177_1_i;
wire na2178_1;
wire na2179_1;
wire na2179_1_i;
wire na2180_1;
wire na2181_1;
wire na2181_1_i;
wire na2182_1;
wire na2183_1;
wire na2183_1_i;
wire na2184_1;
wire na2185_1;
wire na2185_1_i;
wire na2186_1;
wire na2187_1;
wire na2187_1_i;
wire na2188_1;
wire na2189_1;
wire na2189_1_i;
wire na2190_1;
wire na2191_1;
wire na2191_1_i;
wire na2192_1;
wire na2193_1;
wire na2193_1_i;
wire na2194_1;
wire na2195_1;
wire na2195_1_i;
wire na2196_1;
wire na2197_1;
wire na2197_1_i;
wire na2198_1;
wire na2199_1;
wire na2199_1_i;
wire na2200_1;
wire na2201_1;
wire na2201_1_i;
wire na2202_1;
wire na2203_1;
wire na2203_1_i;
wire na2204_1;
wire na2205_1;
wire na2205_1_i;
wire na2206_1;
wire na2207_1;
wire na2207_1_i;
wire na2208_1;
wire na2209_1;
wire na2209_1_i;
wire na2210_1;
wire na2211_1;
wire na2211_1_i;
wire na2212_1;
wire na2213_1;
wire na2213_1_i;
wire na2214_1;
wire na2215_1;
wire na2215_1_i;
wire na2216_1;
wire na2217_1;
wire na2217_1_i;
wire na2218_1;
wire na2219_1;
wire na2219_1_i;
wire na2220_1;
wire na2221_1;
wire na2221_1_i;
wire na2222_1;
wire na2223_1;
wire na2223_1_i;
wire na2224_1;
wire na2225_1;
wire na2225_1_i;
wire na2226_1;
wire na2227_1;
wire na2227_1_i;
wire na2228_1;
wire na2229_1;
wire na2229_1_i;
wire na2230_1;
wire na2231_1;
wire na2231_1_i;
wire na2232_1;
wire na2233_1;
wire na2233_1_i;
wire na2234_1;
wire na2235_1;
wire na2235_1_i;
wire na2236_1;
wire na2237_1;
wire na2237_1_i;
wire na2238_1;
wire na2239_1;
wire na2239_1_i;
wire na2240_1;
wire na2240_1_i;
wire na2241_1;
wire na2242_1;
wire na2242_1_i;
wire na2243_1;
wire na2244_1;
wire na2244_1_i;
wire na2245_1;
wire na2246_1;
wire na2246_1_i;
wire na2248_1;
wire na2249_1;
wire na2250_1;
wire na2251_1;
wire na2251_1_i;
wire na2252_1;
wire na2252_1_i;
wire na2253_1;
wire na2253_1_i;
wire na2254_1;
wire na2254_1_i;
wire na2255_1;
wire na2255_1_i;
wire na2256_1;
wire na2256_1_i;
wire na2257_1;
wire na2262_1;
wire na2263_1;
wire na2264_1;
wire na2265_1;
wire na2266_1;
wire na2267_1;
wire na2268_1;
wire na2269_1;
wire na2270_1;
wire na2271_1;
wire na2272_2;
wire na2273_2;
wire na2274_1;
wire na2275_1;
wire na2276_1;
wire na2277_1;
wire na2278_1;
wire na2279_1;
wire na2280_1;
wire na2281_1;
wire na2282_1;
wire na2283_1;
wire na2284_1;
wire na2285_1;
wire na2286_1;
wire na2287_1;
wire na2288_1;
wire na2289_1;
wire na2290_1;
wire na2291_1;
wire na2292_1;
wire na2293_1;
wire na2294_1;
wire na2295_1;
wire na2296_1;
wire na2297_1;
wire na2298_1;
wire na2299_1;
wire na2300_1;
wire na2301_1;
wire na2302_1;
wire na2303_1;
wire na2306_1;
wire na2309_1;
wire na2309_2;
wire na2310_1;
wire na2311_1;
wire na2312_1;
wire na2314_2;
wire na2315_1;
wire na2316_1;
wire na2316_2;
wire na2317_1;
wire na2318_1;
wire na2318_2;
wire na2320_1;
wire na2321_1;
wire na2321_2;
wire na2322_1;
wire na2322_2;
wire na2324_1;
wire na2325_1;
wire na2327_1;
wire na2327_2;
wire na2328_1;
wire na2331_1;
wire na2332_1;
wire na2332_2;
wire na2333_1;
wire na2334_1;
wire na2335_2;
wire na2336_1;
wire na2337_2;
wire na2338_2;
wire na2339_1;
wire na2340_2;
wire na2341_1;
wire na2342_1;
wire na2344_1;
wire na2344_2;
wire na2346_1;
wire na2348_1;
wire na2348_2;
wire na2349_1;
wire na2351_1;
wire na2351_2;
wire na2352_1;
wire na2354_1;
wire na2354_2;
wire na2355_1;
wire na2357_1;
wire na2357_2;
wire na2358_1;
wire na2360_1;
wire na2361_1;
wire na2361_2;
wire na2362_1;
wire na2363_1;
wire na2364_1;
wire na2364_2;
wire na2366_1;
wire na2367_1;
wire na2369_1;
wire na2369_2;
wire na2370_1;
wire na2372_1;
wire na2372_2;
wire na2373_1;
wire na2376_1;
wire na2378_1;
wire na2378_2;
wire na2379_1;
wire na2380_1;
wire na2383_1;
wire na2383_2;
wire na2384_1;
wire na2385_1;
wire na2386_1;
wire na2388_1;
wire na2389_1;
wire na2390_1;
wire na2390_2;
wire na2391_1;
wire na2392_1;
wire na2393_1;
wire na2394_1;
wire na2395_1;
wire na2396_1;
wire na2397_1;
wire na2398_1;
wire na2399_1;
wire na2400_1;
wire na2401_1;
wire na2402_1;
wire na2403_1;
wire na2404_1;
wire na2405_1;
wire na2406_1;
wire na2407_1;
wire na2408_1;
wire na2409_1;
wire na2410_1;
wire na2411_1;
wire na2412_1;
wire na2413_1;
wire na2414_1;
wire na2415_1;
wire na2416_1;
wire na2417_1;
wire na2418_1;
wire na2419_1;
wire na2420_1;
wire na2421_1;
wire na2422_1;
wire na2422_2;
wire na2423_1;
wire na2423_2;
wire na2424_1;
wire na2424_2;
wire na2425_1;
wire na2425_2;
wire na2426_1;
wire na2426_2;
wire na2427_1;
wire na2427_2;
wire na2428_1;
wire na2428_2;
wire na2429_1;
wire na2429_2;
wire na2430_1;
wire na2430_2;
wire na2431_1;
wire na2431_2;
wire na2432_1;
wire na2432_2;
wire na2433_1;
wire na2433_2;
wire na2434_1;
wire na2434_2;
wire na2435_1;
wire na2435_2;
wire na2436_1;
wire na2436_2;
wire na2437_1;
wire na2437_2;
wire na2438_1;
wire na2438_2;
wire na2439_1;
wire na2439_2;
wire na2440_1;
wire na2440_2;
wire na2441_1;
wire na2441_2;
wire na2442_1;
wire na2442_2;
wire na2443_1;
wire na2443_2;
wire na2444_1;
wire na2444_2;
wire na2445_1;
wire na2445_2;
wire na2446_1;
wire na2446_2;
wire na2447_1;
wire na2447_2;
wire na2448_1;
wire na2448_2;
wire na2449_1;
wire na2449_2;
wire na2450_1;
wire na2450_2;
wire na2451_1;
wire na2451_2;
wire na2454_1;
wire na2455_1;
wire na2456_1;
wire na2456_2;
wire na2457_2;
wire na2459_1;
wire na2460_2;
wire na2462_1;
wire na2463_2;
wire na2465_1;
wire na2466_1;
wire na2468_1;
wire na2469_2;
wire na2471_1;
wire na2472_2;
wire na2474_1;
wire na2475_1;
wire na2477_1;
wire na2478_1;
wire na2479_1;
wire na2480_1;
wire na2481_2;
wire na2482_1;
wire na2484_1;
wire na2486_1;
wire na2488_1;
wire na2490_1;
wire na2492_1;
wire na2494_1;
wire na2496_1;
wire na2498_1;
wire na2500_1;
wire na2502_1;
wire na2504_1;
wire na2506_1;
wire na2508_1;
wire na2510_1;
wire na2512_1;
wire na2514_2;
wire na2515_2;
wire na2516_1;
wire na2517_1;
wire na2518_2;
wire na2519_2;
wire na2520_2;
wire na2520_2_i;
wire na2521_1;
wire na2522_1;
wire na2522_1_i;
wire na2523_1;
wire na2524_1;
wire na2524_1_i;
wire na2525_1;
wire na2526_2;
wire na2526_2_i;
wire na2527_1;
wire na2528_2;
wire na2528_2_i;
wire na2529_1;
wire na2530_1;
wire na2530_1_i;
wire na2531_1;
wire na2532_1;
wire na2532_1_i;
wire na2533_1;
wire na2534_2;
wire na2534_2_i;
wire na2535_1;
wire na2536_1;
wire na2536_1_i;
wire na2537_1;
wire na2537_1_i;
wire na2538_1;
wire na2538_1_i;
wire na2539_1;
wire na2539_1_i;
wire na2540_1;
wire na2540_1_i;
wire na2541_1;
wire na2541_1_i;
wire na2542_1;
wire na2542_1_i;
wire na2543_1;
wire na2543_1_i;
wire na2544_1;
wire na2544_1_i;
wire na2545_2;
wire na2545_2_i;
wire na2546_1;
wire na2546_1_i;
wire na2547_2;
wire na2547_2_i;
wire na2548_1;
wire na2548_1_i;
wire na2549_1;
wire na2549_1_i;
wire na2550_1;
wire na2550_1_i;
wire na2551_2;
wire na2551_2_i;
wire na2552_1;
wire na2552_1_i;
wire na2553_1;
wire na2553_1_i;
wire na2554_1;
wire na2554_1_i;
wire na2555_1;
wire na2555_1_i;
wire na2556_1;
wire na2556_1_i;
wire na2557_1;
wire na2557_1_i;
wire na2558_1;
wire na2558_1_i;
wire na2559_1;
wire na2559_1_i;
wire na2560_1;
wire na2560_1_i;
wire na2561_1;
wire na2561_1_i;
wire na2562_1;
wire na2562_1_i;
wire na2563_1;
wire na2563_1_i;
wire na2564_1;
wire na2564_1_i;
wire na2565_1;
wire na2565_1_i;
wire na2566_1;
wire na2566_1_i;
wire na2567_1;
wire na2567_1_i;
wire na2568_1;
wire na2568_1_i;
wire na2569_1;
wire na2569_1_i;
wire na2570_1;
wire na2570_1_i;
wire na2571_1;
wire na2571_1_i;
wire na2572_1;
wire na2572_1_i;
wire na2573_1;
wire na2573_1_i;
wire na2574_1;
wire na2574_2;
wire na2575_1;
wire na2576_1;
wire na2576_2;
wire na2577_1;
wire na2578_1;
wire na2578_2;
wire na2579_1;
wire na2580_1;
wire na2580_2;
wire na2581_1;
wire na2582_1;
wire na2582_2;
wire na2583_1;
wire na2584_1;
wire na2584_2;
wire na2585_1;
wire na2586_1;
wire na2586_2;
wire na2587_1;
wire na2588_1;
wire na2588_2;
wire na2589_1;
wire na2590_1;
wire na2590_2;
wire na2591_1;
wire na2592_1;
wire na2592_2;
wire na2593_1;
wire na2594_1;
wire na2594_1_i;
wire na2595_1;
wire na2596_1;
wire na2596_1_i;
wire na2597_1;
wire na2597_1_i;
wire na2598_1;
wire na2598_1_i;
wire na2599_1;
wire na2599_1_i;
wire na2600_1;
wire na2600_1_i;
wire na2601_1;
wire na2601_1_i;
wire na2602_1;
wire na2602_1_i;
wire na2603_1;
wire na2603_1_i;
wire na2604_1;
wire na2604_1_i;
wire na2605_1;
wire na2605_1_i;
wire na2606_1;
wire na2606_1_i;
wire na2607_1;
wire na2607_1_i;
wire na2608_1;
wire na2608_1_i;
wire na2609_1;
wire na2609_1_i;
wire na2610_1;
wire na2610_1_i;
wire na2611_1;
wire na2611_1_i;
wire na2612_1;
wire na2612_1_i;
wire na2613_1;
wire na2613_1_i;
wire na2614_1;
wire na2614_1_i;
wire na2615_1;
wire na2615_1_i;
wire na2616_1;
wire na2616_1_i;
wire na2617_1;
wire na2617_1_i;
wire na2618_1;
wire na2618_1_i;
wire na2619_1;
wire na2619_1_i;
wire na2620_1;
wire na2620_1_i;
wire na2621_1;
wire na2621_1_i;
wire na2622_1;
wire na2622_1_i;
wire na2623_1;
wire na2623_1_i;
wire na2624_1;
wire na2624_1_i;
wire na2625_1;
wire na2625_1_i;
wire na2626_1;
wire na2626_1_i;
wire na2627_1;
wire na2627_4;
wire na2659_1;
wire na2659_1_i;
wire na2660_1;
wire na2661_1;
wire na2661_1_i;
wire na2662_1;
wire na2662_1_i;
wire na2663_1;
wire na2664_1;
wire na2664_1_i;
wire na2665_1;
wire na2666_1;
wire na2666_1_i;
wire na2667_1;
wire na2667_1_i;
wire na2668_1;
wire na2668_1_i;
wire na2669_1;
wire na2669_1_i;
wire na2670_1;
wire na2670_1_i;
wire na2671_1;
wire na2671_1_i;
wire na2672_1;
wire na2673_1;
wire na2673_1_i;
wire na2675_1;
wire na2675_1_i;
wire na2676_1;
wire na2677_1;
wire na2677_1_i;
wire na2677_2;
wire na2677_2_i;
wire na2678_1;
wire na2679_2;
wire na2679_2_i;
wire na2680_1;
wire na2681_1;
wire na2681_1_i;
wire na2681_2;
wire na2681_2_i;
wire na2682_1;
wire na2684_1;
wire na2686_1;
wire na2687_1;
wire na2687_1_i;
wire na2687_2;
wire na2687_2_i;
wire na2688_1;
wire na2689_2;
wire na2691_1;
wire na2692_1;
wire na2692_1_i;
wire na2692_2;
wire na2692_2_i;
wire na2693_1;
wire na2693_1_i;
wire na2695_1;
wire na2695_1_i;
wire na2696_2;
wire na2697_1;
wire na2697_1_i;
wire na2698_1;
wire na2698_1_i;
wire na2699_1;
wire na2699_1_i;
wire na2701_1;
wire na2701_1_i;
wire na2702_1;
wire na2702_1_i;
wire na2703_1;
wire na2703_1_i;
wire na2704_1;
wire na2704_1_i;
wire na2705_1;
wire na2705_1_i;
wire na2706_2;
wire na2706_2_i;
wire na2707_1;
wire na2708_1;
wire na2708_1_i;
wire na2709_2;
wire na2710_1;
wire na2710_1_i;
wire na2711_2;
wire na2712_1;
wire na2712_1_i;
wire na2713_1;
wire na2714_1;
wire na2714_1_i;
wire na2715_2;
wire na2716_1;
wire na2716_1_i;
wire na2717_1;
wire na2717_1_i;
wire na2718_1;
wire na2718_1_i;
wire na2718_2;
wire na2718_2_i;
wire na2719_1;
wire na2720_1;
wire na2720_1_i;
wire na2721_1;
wire na2721_1_i;
wire na2722_1;
wire na2723_2;
wire na2723_2_i;
wire na2724_1;
wire na2725_1;
wire na2725_2;
wire na2726_1;
wire na2726_1_i;
wire na2727_1;
wire na2727_1_i;
wire na2728_1;
wire na2728_1_i;
wire na2729_1;
wire na2729_1_i;
wire na2730_1;
wire na2730_1_i;
wire na2731_1;
wire na2731_1_i;
wire na2732_1;
wire na2732_1_i;
wire na2733_1;
wire na2733_1_i;
wire na2734_1;
wire na2734_2;
wire na2735_2;
wire na2735_2_i;
wire na2736_2;
wire na2737_1;
wire na2737_1_i;
wire na2738_1;
wire na2739_1;
wire na2739_1_i;
wire na2740_1;
wire na2740_1_i;
wire na2741_1;
wire na2741_1_i;
wire na2743_1;
wire na2743_1_i;
wire na2744_1;
wire na2744_1_i;
wire na2745_1;
wire na2745_1_i;
wire na2746_2;
wire na2746_2_i;
wire na2747_1;
wire na2748_1;
wire na2748_1_i;
wire na2749_1;
wire na2750_1;
wire na2750_1_i;
wire na2751_1;
wire na2751_2;
wire na2752_1;
wire na2752_1_i;
wire na2753_1;
wire na2753_1_i;
wire na2754_1;
wire na2754_1_i;
wire na2755_1;
wire na2755_1_i;
wire na2756_1;
wire na2756_1_i;
wire na2757_1;
wire na2757_1_i;
wire na2758_1;
wire na2758_1_i;
wire na2759_1;
wire na2759_1_i;
wire na2760_1;
wire na2760_2;
wire na2761_1;
wire na2761_1_i;
wire na2762_1;
wire na2762_1_i;
wire na2763_1;
wire na2764_1;
wire na2764_1_i;
wire na2766_1;
wire na2767_1;
wire na2768_2;
wire na2768_2_i;
wire na2769_2;
wire na2770_1;
wire na2771_1;
wire na2772_2;
wire na2773_1;
wire na2773_1_i;
wire na2774_1;
wire na2774_1_i;
wire na2775_1;
wire na2776_1;
wire na2776_1_i;
wire na2777_2;
wire na2778_1;
wire na2778_1_i;
wire na2779_1;
wire na2780_1;
wire na2780_1_i;
wire na2781_1;
wire na2781_1_i;
wire na2782_1;
wire na2782_1_i;
wire na2783_1;
wire na2783_1_i;
wire na2784_1;
wire na2784_1_i;
wire na2785_1;
wire na2785_1_i;
wire na2786_1;
wire na2786_1_i;
wire na2787_1;
wire na2787_1_i;
wire na2788_1;
wire na2788_1_i;
wire na2789_1;
wire na2789_1_i;
wire na2789_2;
wire na2789_2_i;
wire na2790_1;
wire na2790_1_i;
wire na2791_1;
wire na2791_1_i;
wire na2792_1;
wire na2792_1_i;
wire na2793_1;
wire na2793_1_i;
wire na2794_1;
wire na2794_1_i;
wire na2795_1;
wire na2795_1_i;
wire na2796_1;
wire na2796_1_i;
wire na2797_1;
wire na2797_1_i;
wire na2798_1;
wire na2798_1_i;
wire na2800_1;
wire na2801_1;
wire na2801_1_i;
wire na2802_1;
wire na2802_1_i;
wire na2803_1;
wire na2803_1_i;
wire na2804_1;
wire na2804_1_i;
wire na2805_1;
wire na2805_1_i;
wire na2805_2;
wire na2805_2_i;
wire na2806_1;
wire na2807_2;
wire na2808_2;
wire na2808_2_i;
wire na2809_1;
wire na2810_1;
wire na2811_1;
wire na2811_1_i;
wire na2811_2;
wire na2811_2_i;
wire na2812_1;
wire na2814_1;
wire na2815_1;
wire na2817_1;
wire na2818_1;
wire na2818_1_i;
wire na2818_2;
wire na2818_2_i;
wire na2819_1;
wire na2820_1;
wire na2820_1_i;
wire na2821_1;
wire na2821_1_i;
wire na2822_1;
wire na2823_1;
wire na2823_1_i;
wire na2824_1;
wire na2824_1_i;
wire na2825_1;
wire na2825_1_i;
wire na2826_1;
wire na2826_1_i;
wire na2827_1;
wire na2827_1_i;
wire na2828_1;
wire na2828_1_i;
wire na2829_1;
wire na2829_1_i;
wire na2830_1;
wire na2830_1_i;
wire na2831_2;
wire na2832_1;
wire na2832_1_i;
wire na2833_1;
wire na2833_1_i;
wire na2834_1;
wire na2834_1_i;
wire na2835_1;
wire na2835_1_i;
wire na2835_2;
wire na2835_2_i;
wire na2836_2;
wire na2836_2_i;
wire na2838_1;
wire na2838_1_i;
wire na2839_1;
wire na2840_1;
wire na2841_2;
wire na2842_2;
wire na2843_1;
wire na2844_2;
wire na2845_2;
wire na2846_2;
wire na2847_1;
wire na2848_2;
wire na2849_1;
wire na2850_2;
wire na2851_2;
wire na2852_1;
wire na2853_1;
wire na2854_2;
wire na2855_2;
wire na2856_1;
wire na2857_2;
wire na2858_1;
wire na2859_1;
wire na2860_2;
wire na2861_1;
wire na2862_1;
wire na2863_2;
wire na2864_2;
wire na2865_2;
wire na2866_1;
wire na2867_2;
wire na2868_1;
wire na2869_1;
wire na2870_2;
wire na2871_2;
wire na2872_1;
wire na2873_1;
wire na2874_2;
wire na2875_1;
wire na2876_2;
wire na2877_2;
wire na2878_2;
wire na2879_1;
wire na2880_2;
wire na2881_1;
wire na2882_2;
wire na2883_1;
wire na2884_2;
wire na2885_1;
wire na2886_2;
wire na2887_1;
wire na2888_2;
wire na2889_1;
wire na2890_1;
wire na2891_2;
wire na2892_2;
wire na2894_2;
wire na2894_2_i;
wire na2895_1;
wire na2895_1_i;
wire na2897_1;
wire na2897_1_i;
wire na2897_2;
wire na2897_2_i;
wire na2898_1;
wire na2898_1_i;
wire na2898_2;
wire na2898_2_i;
wire na2899_1;
wire na2899_1_i;
wire na2899_2;
wire na2899_2_i;
wire na2900_1;
wire na2900_1_i;
wire na2900_2;
wire na2900_2_i;
wire na2901_1;
wire na2901_1_i;
wire na2901_2;
wire na2901_2_i;
wire na2902_1;
wire na2902_1_i;
wire na2904_1;
wire na2904_1_i;
wire na2904_2;
wire na2904_2_i;
wire na2906_1;
wire na2906_1_i;
wire na2907_1;
wire na2907_1_i;
wire na2907_2;
wire na2907_2_i;
wire na2908_1;
wire na2908_1_i;
wire na2909_1;
wire na2909_1_i;
wire na2910_1;
wire na2910_1_i;
wire na2911_1;
wire na2911_1_i;
wire na2912_1;
wire na2912_1_i;
wire na2913_1;
wire na2913_1_i;
wire na2914_1;
wire na2914_1_i;
wire na2915_1;
wire na2915_1_i;
wire na2917_2;
wire na2917_2_i;
wire na2918_1;
wire na2918_1_i;
wire na2919_1;
wire na2919_1_i;
wire na2920_2;
wire na2920_2_i;
wire na2921_1;
wire na2922_1;
wire na2922_1_i;
wire na2923_1;
wire na2924_1;
wire na2924_1_i;
wire na2925_1;
wire na2925_1_i;
wire na2926_1;
wire na2926_1_i;
wire na2927_1;
wire na2927_1_i;
wire na2928_1;
wire na2928_1_i;
wire na2929_1;
wire na2929_1_i;
wire na2930_1;
wire na2930_1_i;
wire na2931_1;
wire na2931_1_i;
wire na2932_1;
wire na2933_2;
wire na2933_2_i;
wire na2935_1;
wire na2935_1_i;
wire na2936_1;
wire na2936_1_i;
wire na2937_2;
wire na2937_2_i;
wire na2938_1;
wire na2938_1_i;
wire na2939_1;
wire na2939_1_i;
wire na2940_1;
wire na2940_1_i;
wire na2941_1;
wire na2941_1_i;
wire na2942_1;
wire na2942_1_i;
wire na2943_1;
wire na2943_1_i;
wire na2944_1;
wire na2944_1_i;
wire na2945_1;
wire na2945_1_i;
wire na2946_1;
wire na2946_1_i;
wire na2947_1;
wire na2947_1_i;
wire na2948_2;
wire na2948_2_i;
wire na2949_1;
wire na2950_1;
wire na2950_1_i;
wire na2951_2;
wire na2951_2_i;
wire na2952_2;
wire na2953_1;
wire na2953_1_i;
wire na2953_2;
wire na2953_2_i;
wire na2954_2;
wire na2955_1;
wire na2955_1_i;
wire na2956_1;
wire na2956_1_i;
wire na2957_1;
wire na2957_1_i;
wire na2959_2;
wire na2960_1;
wire na2960_1_i;
wire na2961_1;
wire na2962_1;
wire na2962_1_i;
wire na2963_1;
wire na2963_1_i;
wire na2964_1;
wire na2964_1_i;
wire na2965_1;
wire na2965_1_i;
wire na2966_1;
wire na2966_1_i;
wire na2967_1;
wire na2967_1_i;
wire na2968_1;
wire na2968_1_i;
wire na2969_1;
wire na2969_1_i;
wire na2970_1;
wire na2970_1_i;
wire na2971_1;
wire na2971_1_i;
wire na2972_1;
wire na2972_1_i;
wire na2972_2;
wire na2972_2_i;
wire na2973_1;
wire na2974_1;
wire na2974_1_i;
wire na2975_1;
wire na2975_1_i;
wire na2976_1;
wire na2976_1_i;
wire na2977_1;
wire na2977_1_i;
wire na2978_1;
wire na2978_1_i;
wire na2979_1;
wire na2979_1_i;
wire na2980_2;
wire na2980_2_i;
wire na2981_1;
wire na2981_1_i;
wire na2982_2;
wire na2983_1;
wire na2983_1_i;
wire na2984_1;
wire na2986_1;
wire na2986_2;
wire na2987_1;
wire na2987_1_i;
wire na2989_1;
wire na2989_1_i;
wire na2990_2;
wire na2991_1;
wire na2991_1_i;
wire na2992_1;
wire na2992_1_i;
wire na2993_1;
wire na2993_1_i;
wire na2994_1;
wire na2994_1_i;
wire na2995_1;
wire na2995_1_i;
wire na2996_1;
wire na2996_1_i;
wire na2998_1;
wire na3000_1;
wire na3001_1;
wire na3001_1_i;
wire na3002_1;
wire na3002_1_i;
wire na3003_1;
wire na3003_1_i;
wire na3003_2;
wire na3003_2_i;
wire na3006_1;
wire na3006_1_i;
wire na3006_2;
wire na3006_2_i;
wire na3008_1;
wire na3008_1_i;
wire na3009_1;
wire na3009_1_i;
wire na3010_1;
wire na3010_1_i;
wire na3011_1;
wire na3011_1_i;
wire na3012_1;
wire na3012_1_i;
wire na3013_2;
wire na3013_2_i;
wire na3014_2;
wire na3014_2_i;
wire na3015_1;
wire na3016_1;
wire na3016_1_i;
wire na3017_1;
wire na3017_1_i;
wire na3018_1;
wire na3018_1_i;
wire na3018_2;
wire na3018_2_i;
wire na3020_1;
wire na3020_1_i;
wire na3020_2;
wire na3020_2_i;
wire na3022_1;
wire na3022_1_i;
wire na3022_2;
wire na3022_2_i;
wire na3024_1;
wire na3024_1_i;
wire na3024_2;
wire na3024_2_i;
wire na3026_1;
wire na3026_1_i;
wire na3026_2;
wire na3026_2_i;
wire na3027_1;
wire na3027_1_i;
wire na3029_2;
wire na3029_2_i;
wire na3031_1;
wire na3031_1_i;
wire na3031_2;
wire na3031_2_i;
wire na3032_1;
wire na3032_1_i;
wire na3032_2;
wire na3032_2_i;
wire na3034_1;
wire na3034_1_i;
wire na3035_1;
wire na3036_1;
wire na3036_1_i;
wire na3037_1;
wire na3038_1;
wire na3038_1_i;
wire na3039_1;
wire na3040_1;
wire na3040_1_i;
wire na3041_1;
wire na3042_1;
wire na3042_1_i;
wire na3043_1;
wire na3044_1;
wire na3044_1_i;
wire na3045_1;
wire na3046_1;
wire na3046_1_i;
wire na3047_1;
wire na3048_1;
wire na3048_1_i;
wire na3049_1;
wire na3050_1;
wire na3050_1_i;
wire na3051_1;
wire na3052_1;
wire na3052_1_i;
wire na3053_1;
wire na3054_1;
wire na3054_1_i;
wire na3055_1;
wire na3056_1;
wire na3056_1_i;
wire na3057_1;
wire na3058_1;
wire na3058_1_i;
wire na3059_1;
wire na3060_1;
wire na3060_1_i;
wire na3061_1;
wire na3062_1;
wire na3062_1_i;
wire na3063_1;
wire na3064_1;
wire na3064_1_i;
wire na3064_2;
wire na3064_2_i;
wire na3065_1;
wire na3065_1_i;
wire na3066_1;
wire na3066_1_i;
wire na3068_1;
wire na3068_1_i;
wire na3069_1;
wire na3070_1;
wire na3070_1_i;
wire na3071_1;
wire na3071_1_i;
wire na3072_1;
wire na3072_1_i;
wire na3073_1;
wire na3073_1_i;
wire na3074_1;
wire na3074_1_i;
wire na3075_1;
wire na3075_1_i;
wire na3076_1;
wire na3076_1_i;
wire na3077_1;
wire na3077_1_i;
wire na3078_1;
wire na3079_1;
wire na3079_1_i;
wire na3080_1;
wire na3081_1;
wire na3081_1_i;
wire na3082_1;
wire na3083_1;
wire na3083_1_i;
wire na3084_1;
wire na3085_1;
wire na3085_1_i;
wire na3086_1;
wire na3087_1;
wire na3087_1_i;
wire na3088_1;
wire na3089_1;
wire na3089_1_i;
wire na3090_1;
wire na3091_1;
wire na3091_1_i;
wire na3092_1;
wire na3093_1;
wire na3093_1_i;
wire na3094_1;
wire na3095_1;
wire na3095_1_i;
wire na3096_1;
wire na3097_1;
wire na3097_1_i;
wire na3098_1;
wire na3099_1;
wire na3099_1_i;
wire na3100_1;
wire na3101_1;
wire na3101_1_i;
wire na3102_1;
wire na3103_1;
wire na3103_1_i;
wire na3104_1;
wire na3105_1;
wire na3105_1_i;
wire na3106_1;
wire na3107_1;
wire na3107_1_i;
wire na3107_2;
wire na3107_2_i;
wire na3108_2;
wire na3109_1;
wire na3109_1_i;
wire na3110_1;
wire na3110_1_i;
wire na3111_1;
wire na3111_1_i;
wire na3112_1;
wire na3112_1_i;
wire na3113_1;
wire na3113_1_i;
wire na3114_1;
wire na3114_1_i;
wire na3115_1;
wire na3115_1_i;
wire na3115_2;
wire na3115_2_i;
wire na3116_1;
wire na3116_1_i;
wire na3117_1;
wire na3117_1_i;
wire na3118_1;
wire na3118_1_i;
wire na3119_1;
wire na3119_1_i;
wire na3121_1;
wire na3121_1_i;
wire na3122_1;
wire na3122_1_i;
wire na3122_2;
wire na3122_2_i;
wire na3123_1;
wire na3123_1_i;
wire na3124_1;
wire na3124_1_i;
wire na3125_1;
wire na3125_1_i;
wire na3126_1;
wire na3126_1_i;
wire na3127_1;
wire na3127_1_i;
wire na3127_2;
wire na3127_2_i;
wire na3128_1;
wire na3128_1_i;
wire na3129_1;
wire na3129_1_i;
wire na3130_1;
wire na3130_1_i;
wire na3131_1;
wire na3131_1_i;
wire na3131_2;
wire na3131_2_i;
wire na3132_1;
wire na3132_1_i;
wire na3134_1;
wire na3134_1_i;
wire na3136_1;
wire na3136_1_i;
wire na3137_1;
wire na3137_1_i;
wire na3137_2;
wire na3137_2_i;
wire na3138_1;
wire na3138_1_i;
wire na3139_1;
wire na3139_1_i;
wire na3140_1;
wire na3140_1_i;
wire na3141_1;
wire na3141_1_i;
wire na3142_2;
wire na3142_2_i;
wire na3143_1;
wire na3143_1_i;
wire na3145_1;
wire na3145_1_i;
wire na3146_1;
wire na3146_1_i;
wire na3147_1;
wire na3147_1_i;
wire na3148_1;
wire na3148_1_i;
wire na3149_1;
wire na3149_1_i;
wire na3150_1;
wire na3150_1_i;
wire na3151_1;
wire na3151_1_i;
wire na3152_1;
wire na3152_1_i;
wire na3153_1;
wire na3153_1_i;
wire na3154_1;
wire na3154_1_i;
wire na3155_1;
wire na3155_1_i;
wire na3156_1;
wire na3156_1_i;
wire na3158_1;
wire na3158_1_i;
wire na3159_1;
wire na3159_1_i;
wire na3159_2;
wire na3159_2_i;
wire na3161_1;
wire na3161_1_i;
wire na3162_1;
wire na3162_1_i;
wire na3162_2;
wire na3162_2_i;
wire na3163_1;
wire na3163_1_i;
wire na3164_1;
wire na3164_1_i;
wire na3165_1;
wire na3165_1_i;
wire na3166_1;
wire na3166_1_i;
wire na3167_1;
wire na3167_1_i;
wire na3168_1;
wire na3168_1_i;
wire na3169_1;
wire na3169_1_i;
wire na3170_1;
wire na3170_1_i;
wire na3171_1;
wire na3171_1_i;
wire na3172_1;
wire na3172_1_i;
wire na3173_1;
wire na3173_1_i;
wire na3173_2;
wire na3173_2_i;
wire na3174_1;
wire na3174_1_i;
wire na3175_1;
wire na3175_1_i;
wire na3177_1;
wire na3177_1_i;
wire na3178_2;
wire na3178_2_i;
wire na3179_1;
wire na3180_1;
wire na3180_1_i;
wire na3181_2;
wire na3182_1;
wire na3182_1_i;
wire na3182_2;
wire na3182_2_i;
wire na3183_1;
wire na3183_1_i;
wire na3185_1;
wire na3185_1_i;
wire na3186_2;
wire na3186_2_i;
wire na3187_1;
wire na3188_1;
wire na3188_1_i;
wire na3188_2;
wire na3188_2_i;
wire na3189_1;
wire na3189_1_i;
wire na3190_1;
wire na3190_1_i;
wire na3191_1;
wire na3191_1_i;
wire na3192_1;
wire na3192_1_i;
wire na3193_1;
wire na3193_1_i;
wire na3194_1;
wire na3194_1_i;
wire na3195_1;
wire na3195_1_i;
wire na3196_1;
wire na3196_1_i;
wire na3197_1;
wire na3197_1_i;
wire na3198_1;
wire na3198_1_i;
wire na3200_1;
wire na3200_1_i;
wire na3201_1;
wire na3201_1_i;
wire na3203_1;
wire na3203_1_i;
wire na3204_1;
wire na3204_1_i;
wire na3205_1;
wire na3205_1_i;
wire na3207_1;
wire na3207_1_i;
wire na3208_1;
wire na3208_1_i;
wire na3210_1;
wire na3210_1_i;
wire na3211_1;
wire na3211_1_i;
wire na3212_1;
wire na3212_1_i;
wire na3213_1;
wire na3214_1;
wire na3214_2;
wire na3215_1;
wire na3216_2;
wire na3216_2_i;
wire na3217_1;
wire na3218_2;
wire na3219_1;
wire na3219_1_i;
wire na3219_2;
wire na3219_2_i;
wire na3220_1;
wire na3222_1;
wire na3222_1_i;
wire na3224_2;
wire na3225_1;
wire na3226_1;
wire na3226_2;
wire na3227_2;
wire na3227_2_i;
wire na3228_1;
wire na3229_2;
wire na3230_2;
wire na3231_1;
wire na3232_1;
wire na3233_2;
wire na3234_2;
wire na3237_1;
wire na3238_2;
wire na3239_1;
wire na3240_2;
wire na3241_1;
wire na3242_1;
wire na3243_1;
wire na3244_2;
wire na3247_1;
wire na3248_2;
wire na3249_2;
wire na3250_1;
wire na3251_2;
wire na3253_1;
wire na3254_2;
wire na3255_1;
wire na3256_1;
wire na3256_1_i;
wire na3257_1;
wire na3258_1;
wire na3258_2;
wire na3259_1;
wire na3259_1_i;
wire na3262_1;
wire na3262_1_i;
wire na3263_1;
wire na3263_1_i;
wire na3264_1;
wire na3264_1_i;
wire na3265_1;
wire na3265_1_i;
wire na3266_1;
wire na3266_1_i;
wire na3268_2;
wire na3268_2_i;
wire na3269_2;
wire na3269_2_i;
wire na3270_1;
wire na3270_1_i;
wire na3272_2;
wire na3273_1;
wire na3274_2;
wire na3275_1;
wire na3276_1;
wire na3276_1_i;
wire na3277_1;
wire na3278_2;
wire na3279_1;
wire na3280_1;
wire na3281_1;
wire na3282_1;
wire na3283_1;
wire na3284_2;
wire na3285_1;
wire na3286_1;
wire na3287_2;
wire na3288_1;
wire na3289_2;
wire na3290_1;
wire na3290_1_i;
wire na3292_1;
wire na3292_1_i;
wire na3296_1;
wire na3297_1;
wire na3297_1_i;
wire na3297_2;
wire na3297_2_i;
wire na3298_1;
wire na3299_2;
wire na3299_2_i;
wire na3300_2;
wire na3301_1;
wire na3301_1_i;
wire na3302_1;
wire na3303_1;
wire na3304_2;
wire na3305_1;
wire na3305_1_i;
wire na3307_1;
wire na3307_2;
wire na3308_1;
wire na3308_1_i;
wire na3309_1;
wire na3309_1_i;
wire na3309_2;
wire na3309_2_i;
wire na3311_1;
wire na3313_1;
wire na3313_1_i;
wire na3313_2;
wire na3313_2_i;
wire na3315_1;
wire na3315_1_i;
wire na3316_1;
wire na3317_1;
wire na3317_1_i;
wire na3319_1;
wire na3319_1_i;
wire na3321_1;
wire na3321_1_i;
wire na3323_1;
wire na3323_1_i;
wire na3324_1;
wire na3324_1_i;
wire na3325_1;
wire na3325_1_i;
wire na3326_2;
wire na3326_2_i;
wire na3327_2;
wire na3327_2_i;
wire na3328_1;
wire na3328_1_i;
wire na3329_2;
wire na3329_2_i;
wire na3330_1;
wire na3330_1_i;
wire na3331_1;
wire na3332_1;
wire na3333_1;
wire na3333_2;
wire na3334_2;
wire na3335_2;
wire na3337_1;
wire na3339_2;
wire na3340_1;
wire na3341_1;
wire na3342_1;
wire na3343_1;
wire na3343_1_i;
wire na3345_1;
wire na3345_1_i;
wire na3347_2;
wire na3348_1;
wire na3349_2;
wire na3350_1;
wire na3351_2;
wire na3352_2;
wire na3352_2_i;
wire na3353_1;
wire na3354_1;
wire na3354_1_i;
wire na3356_1;
wire na3356_1_i;
wire na3357_1;
wire na3357_1_i;
wire na3359_2;
wire na3360_1;
wire na3361_1;
wire na3362_1;
wire na3363_1;
wire na3364_1;
wire na3365_2;
wire na3366_1;
wire na3367_1;
wire na3368_1;
wire na3369_2;
wire na3370_1;
wire na3371_2;
wire na3372_1;
wire na3373_1;
wire na3374_1;
wire na3375_2;
wire na3376_1;
wire na3377_1;
wire na3378_1;
wire na3379_2;
wire na3380_1;
wire na3381_2;
wire na3382_1;
wire na3383_1;
wire na3384_1;
wire na3385_2;
wire na3386_1;
wire na3387_1;
wire na3388_1;
wire na3389_1;
wire na3390_1;
wire na3391_2;
wire na3392_1;
wire na3393_1;
wire na3394_1;
wire na3395_1;
wire na3396_1;
wire na3397_1;
wire na3398_1;
wire na3399_1;
wire na3400_1;
wire na3401_1;
wire na3402_1;
wire na3403_2;
wire na3404_1;
wire na3405_1;
wire na3406_1;
wire na3407_2;
wire na3408_1;
wire na3409_2;
wire na3410_1;
wire na3411_1;
wire na3412_1;
wire na3413_2;
wire na3414_1;
wire na3415_1;
wire na3416_1;
wire na3417_2;
wire na3418_1;
wire na3419_2;
wire na3420_1;
wire na3421_1;
wire na3423_1;
wire na3423_1_i;
wire na3424_2;
wire na3424_2_i;
wire na3486_1;
wire na3487_1;
wire na3488_1;
wire na3489_1;
wire na3490_1;
wire na3491_1;
wire na3492_1;
wire na3494_1;
wire na3494_2;
wire na3496_1;
wire na3496_2;
wire na3497_1;
wire na3498_1;
wire na3499_1;
wire na3499_2;
wire na3501_1;
wire na3503_1;
wire na3504_1;
wire na3508_1;
wire na3512_1;
wire na3514_1;
wire na3521_1;
wire na3525_1;
wire na3526_1;
wire na3527_1;
wire na3529_1;
wire na3530_1;
wire na3531_1;
wire na3532_1;
wire na3535_1;
wire na3537_1;
wire na3539_1;
wire na3540_1;
wire na3542_1;
wire na3543_1;
wire na3544_1;
wire na3546_1;
wire na3547_1;
wire na3548_1;
wire na3548_1_i;
wire na3549_1;
wire na3550_1;
wire na3552_2;
wire na3554_1;
wire na3554_1_i;
wire na3555_1;
wire na3559_1;
wire na3559_1_i;
wire na3560_2;
wire na3561_1;
wire na3562_1;
wire na3562_1_i;
wire na3563_1;
wire na3564_1;
wire na3565_1;
wire na3566_1;
wire na3567_1;
wire na3568_1;
wire na3569_1;
wire na3570_1;
wire na3571_1;
wire na3572_1;
wire na3573_1;
wire na3574_1;
wire na3575_1;
wire na3576_1;
wire na3577_1;
wire na3578_1;
wire na3579_1;
wire na3580_1;
wire na3581_1;
wire na3582_1;
wire na3583_1;
wire na3584_1;
wire na3585_1;
wire na3586_2;
wire na3587_1;
wire na3588_1;
wire na3588_1_i;
wire na3588_2;
wire na3588_2_i;
wire na3589_2;
wire na3590_2;
wire na3590_2_i;
wire na3592_1;
wire na3593_2;
wire na3594_1;
wire na3594_1_i;
wire na3595_1;
wire na3596_2;
wire na3596_2_i;
wire na3597_1;
wire na3598_2;
wire na3598_2_i;
wire na3599_2;
wire na3600_1;
wire na3600_1_i;
wire na3603_1;
wire na3605_1;
wire na3607_1;
wire na3608_1;
wire na3609_1;
wire na3610_2;
wire na3611_1;
wire na3612_1;
wire na3613_4;
wire na3615_4;
wire na3617_4;
wire na3618_4;
wire na3619_1;
wire na3619_4;
wire na3620_1;
wire na3620_4;
wire na3621_1;
wire na3640_4;
wire na3644_4;
wire na3646_1;
wire na3651_4;
wire na3653_4;
wire na3655_4;
wire na3657_4;
wire na3659_4;
wire na3660_4;
wire na3661_1;
wire na3661_4;
wire na3662_1;
wire na3662_4;
wire na3663_1;
wire na3663_4;
wire na3664_1;
wire na3665_1;
wire na3682_4;
wire na3686_4;
wire na3688_1;
wire na3693_4;
wire na3695_4;
wire na3697_1;
wire na3697_4;
wire na3698_1;
wire na3698_2;
wire na3698_4;
wire na3700_1;
wire na3701_1;
wire na3701_4;
wire na3703_1;
wire na3703_2;
wire na3703_4;
wire na3705_1;
wire na3705_2;
wire na3705_4;
wire na3707_1;
wire na3707_2;
wire na3707_4;
wire na3709_1;
wire na3709_2;
wire na3709_4;
wire na3711_1;
wire na3711_2;
wire na3711_4;
wire na3712_1;
wire na3712_2;
wire na3712_4;
wire na3714_1;
wire na3714_2;
wire na3714_4;
wire na3716_1;
wire na3716_2;
wire na3716_4;
wire na3718_1;
wire na3718_2;
wire na3718_4;
wire na3720_1;
wire na3720_2;
wire na3720_4;
wire na3722_1;
wire na3722_4;
wire na3724_1;
wire na3724_4;
wire na3725_1;
wire na3725_2;
wire na3725_4;
wire na3727_1;
wire na3727_2;
wire na3727_4;
wire na3729_1;
wire na3729_2;
wire na3729_4;
wire na3731_1;
wire na3731_2;
wire na3731_4;
wire na3732_1;
wire na3733_1;
wire na3733_2;
wire na3733_4;
wire na3735_1;
wire na3735_2;
wire na3735_4;
wire na3737_1;
wire na3737_2;
wire na3737_4;
wire na3739_1;
wire na3740_1;
wire na3740_4;
wire na3742_1;
wire na3742_2;
wire na3742_4;
wire na3744_1;
wire na3744_2;
wire na3744_4;
wire na3746_1;
wire na3746_2;
wire na3746_4;
wire na3748_1;
wire na3748_2;
wire na3748_4;
wire na3750_1;
wire na3750_2;
wire na3750_4;
wire na3751_1;
wire na3751_2;
wire na3751_4;
wire na3753_1;
wire na3753_2;
wire na3753_4;
wire na3755_1;
wire na3755_2;
wire na3755_4;
wire na3757_1;
wire na3757_2;
wire na3757_4;
wire na3759_1;
wire na3759_2;
wire na3759_4;
wire na3761_1;
wire na3761_2;
wire na3761_4;
wire na3764_1;
wire na3765_1;
wire na3765_2;
wire na3765_4;
wire na3767_1;
wire na3767_2;
wire na3767_4;
wire na3769_1;
wire na3769_2;
wire na3769_4;
wire na3771_1;
wire na3771_2;
wire na3771_4;
wire na3772_1;
wire na3772_4;
wire na3774_1;
wire na3774_2;
wire na3774_4;
wire na3776_1;
wire na3776_2;
wire na3776_4;
wire na3778_1;
wire na3778_2;
wire na3778_4;
wire na3780_1;
wire na3780_2;
wire na3780_4;
wire na3782_1;
wire na3782_2;
wire na3782_4;
wire na3783_1;
wire na3783_2;
wire na3783_4;
wire na3785_1;
wire na3785_2;
wire na3785_4;
wire na3787_1;
wire na3787_2;
wire na3787_4;
wire na3789_1;
wire na3789_2;
wire na3789_4;
wire na3791_1;
wire na3791_2;
wire na3791_4;
wire na3793_1;
wire na3793_2;
wire na3793_4;
wire na3796_1;
wire na3796_4;
wire na3797_1;
wire na3797_4;
wire na3798_1;
wire na3798_2;
wire na3798_4;
wire na3800_1;
wire na3800_2;
wire na3800_4;
wire na3802_1;
wire na3802_2;
wire na3802_4;
wire na3804_1;
wire na3804_2;
wire na3804_4;
wire na3805_1;
wire na3807_1;
wire na3807_2;
wire na3807_4;
wire na3809_1;
wire na3809_2;
wire na3809_4;
wire na3811_1;
wire na3811_2;
wire na3811_4;
wire na3813_1;
wire na3813_2;
wire na3813_4;
wire na3815_1;
wire na3815_2;
wire na3815_4;
wire na3816_1;
wire na3816_2;
wire na3816_4;
wire na3818_1;
wire na3818_2;
wire na3818_4;
wire na3820_1;
wire na3820_2;
wire na3820_4;
wire na3822_1;
wire na3822_2;
wire na3822_4;
wire na3824_1;
wire na3824_2;
wire na3824_4;
wire na3826_1;
wire na3826_2;
wire na3826_4;
wire na3829_1;
wire na3829_4;
wire na3830_1;
wire na3830_4;
wire na3831_1;
wire na3831_2;
wire na3831_4;
wire na3833_1;
wire na3833_2;
wire na3833_4;
wire na3835_1;
wire na3835_2;
wire na3835_4;
wire na3837_1;
wire na3837_2;
wire na3837_4;
wire na3838_1;
wire na3839_1;
wire na3839_2;
wire na3839_4;
wire na3841_1;
wire na3842_1;
wire na3842_4;
wire na3843_1;
wire na3843_2;
wire na3843_4;
wire na3845_1;
wire na3846_1;
wire na3846_4;
wire na3847_1;
wire na3847_2;
wire na3847_4;
wire na3849_1;
wire na3849_2;
wire na3851_1;
wire na3851_4;
wire na3852_1;
wire na3852_2;
wire na3852_4;
wire na3854_1;
wire na3855_1;
wire na3855_4;
wire na3856_1;
wire na3856_2;
wire na3856_4;
wire na3858_1;
wire na3859_1;
wire na3859_4;
wire na3860_1;
wire na3860_2;
wire na3860_4;
wire na3862_1;
wire na3862_2;
wire na3864_1;
wire na3864_4;
wire na3865_1;
wire na3865_2;
wire na3867_1;
wire na3867_4;
wire na3868_1;
wire na3868_2;
wire na3870_1;
wire na3870_4;
wire na3871_1;
wire na3871_2;
wire na3873_1;
wire na3873_4;
wire na3874_1;
wire na3874_2;
wire na3874_4;
wire na3876_1;
wire na3877_1;
wire na3877_4;
wire na3878_1;
wire na3878_2;
wire na3880_1;
wire na3880_4;
wire na3881_1;
wire na3881_2;
wire na3881_4;
wire na3883_1;
wire na3884_1;
wire na3884_4;
wire na3885_1;
wire na3885_2;
wire na3887_1;
wire na3887_4;
wire na3888_1;
wire na3888_2;
wire na3888_4;
wire na3890_1;
wire na3891_1;
wire na3891_4;
wire na3892_1;
wire na3892_2;
wire na3892_4;
wire na3894_1;
wire na3895_1;
wire na3895_4;
wire na3896_1;
wire na3896_2;
wire na3898_1;
wire na3898_4;
wire na3899_1;
wire na3899_2;
wire na3899_4;
wire na3901_1;
wire na3902_1;
wire na3902_4;
wire na3903_1;
wire na3903_2;
wire na3905_1;
wire na3905_4;
wire na3906_1;
wire na3906_2;
wire na3906_4;
wire na3908_1;
wire na3909_1;
wire na3909_2;
wire na3909_4;
wire na3910_1;
wire na3910_2;
wire na3910_4;
wire na3912_1;
wire na3912_2;
wire na3912_4;
wire na3914_1;
wire na3914_2;
wire na3914_4;
wire na3916_1;
wire na3916_2;
wire na3916_4;
wire na3918_1;
wire na3918_2;
wire na3918_4;
wire na3921_1;
wire na3921_2;
wire na3921_4;
wire na3923_1;
wire na3923_2;
wire na3923_4;
wire na3925_1;
wire na3925_2;
wire na3925_4;
wire na3927_1;
wire na3927_2;
wire na3927_4;
wire na3929_1;
wire na3929_2;
wire na3931_1;
wire na3931_2;
wire na3931_4;
wire na3933_1;
wire na3933_2;
wire na3933_4;
wire na3935_1;
wire na3935_2;
wire na3935_4;
wire na3937_1;
wire na3937_2;
wire na3937_4;
wire na3939_4;
wire na3941_1;
wire na3941_1_i;
wire na3941_2;
wire na3941_4;
wire na3943_1;
wire na3943_1_i;
wire na3943_2;
wire na3943_4;
wire na3945_1;
wire na3945_1_i;
wire na3945_2;
wire na3945_4;
wire na3947_1;
wire na3947_1_i;
wire na3947_2;
wire na3947_4;
wire na3949_1;
wire na3949_1_i;
wire na3949_2;
wire na3949_4;
wire na3950_1;
wire na3950_1_i;
wire na3950_4;
wire na3952_1;
wire na3952_1_i;
wire na3952_2;
wire na3952_4;
wire na3954_1;
wire na3954_1_i;
wire na3954_2;
wire na3954_4;
wire na3956_1;
wire na3956_1_i;
wire na3956_2;
wire na3956_4;
wire na3958_1;
wire na3958_1_i;
wire na3958_2;
wire na3958_4;
wire na3960_1;
wire na3960_1_i;
wire na3960_2;
wire na3960_4;
wire na3961_1;
wire na3961_1_i;
wire na3961_4;
wire na3963_1;
wire na3963_1_i;
wire na3964_1;
wire na3964_1_i;
wire na3964_4;
wire na3965_1;
wire na3965_1_i;
wire na3965_4;
wire na3966_1;
wire na3966_1_i;
wire na3966_2;
wire na3966_4;
wire na3968_1;
wire na3968_1_i;
wire na3968_2;
wire na3968_4;
wire na3970_1;
wire na3970_1_i;
wire na3970_2;
wire na3970_4;
wire na3971_1;
wire na3971_4;
wire na3972_1;
wire na3972_2;
wire na3974_1;
wire na3974_4;
wire na3975_1;
wire na3975_2;
wire na3977_1;
wire na3977_2;
wire na3977_4;
wire na3979_1;
wire na3980_1;
wire na3980_2;
wire na3980_4;
wire na3982_1;
wire na3983_1;
wire na3983_4;
wire na3984_1;
wire na3984_1_i;
wire na3984_2;
wire na3984_4;
wire na3986_1;
wire na3986_1_i;
wire na3986_2;
wire na3988_1;
wire na3988_4;
wire na3990_1;
wire na3990_2;
wire na3990_4;
wire na3992_1;
wire na3992_2;
wire na3992_4;
wire na3994_1;
wire na3994_2;
wire na3994_4;
wire na3996_1;
wire na3996_2;
wire na3996_4;
wire na3998_1;
wire na3998_2;
wire na3998_4;
wire na3999_1;
wire na3999_2;
wire na3999_4;
wire na4001_1;
wire na4001_2;
wire na4001_4;
wire na4003_1;
wire na4003_2;
wire na4003_4;
wire na4005_1;
wire na4005_2;
wire na4005_4;
wire na4007_1;
wire na4007_2;
wire na4007_4;
wire na4009_1;
wire na4009_2;
wire na4009_4;
wire na4012_1;
wire na4013_1;
wire na4013_2;
wire na4013_4;
wire na4015_1;
wire na4015_2;
wire na4015_4;
wire na4017_1;
wire na4017_2;
wire na4017_4;
wire na4019_1;
wire na4019_2;
wire na4019_4;
wire na4020_1;
wire na4020_4;
wire na4021_1;
wire na4021_2;
wire na4021_4;
wire na4023_1;
wire na4023_2;
wire na4025_1;
wire na4025_4;
wire na4026_1;
wire na4026_4;
wire na4027_1;
wire na4027_4;
wire na4028_1;
wire na4028_4;
wire na4029_1;
wire na4029_4;
wire na4030_1;
wire na4030_4;
wire na4031_1;
wire na4031_4;
wire na4033_1;
wire na4033_2;
wire na4033_4;
wire na4035_1;
wire na4035_2;
wire na4035_4;
wire na4037_1;
wire na4037_2;
wire na4037_4;
wire na4039_1;
wire na4039_2;
wire na4039_4;
wire na4041_1;
wire na4041_2;
wire na4041_4;
wire na4042_1;
wire na4042_2;
wire na4042_4;
wire na4044_1;
wire na4044_2;
wire na4044_4;
wire na4046_1;
wire na4046_2;
wire na4046_4;
wire na4048_1;
wire na4048_2;
wire na4048_4;
wire na4050_1;
wire na4050_2;
wire na4050_4;
wire na4052_1;
wire na4052_2;
wire na4052_4;
wire na4055_1;
wire na4056_1;
wire na4056_2;
wire na4056_4;
wire na4058_1;
wire na4058_2;
wire na4058_4;
wire na4060_1;
wire na4060_2;
wire na4060_4;
wire na4062_1;
wire na4062_2;
wire na4062_4;
wire na4063_1;
wire na4063_4;
wire na4064_1;
wire na4064_2;
wire na4064_4;
wire na4066_1;
wire na4066_2;
wire na4068_1;
wire na4068_4;
wire na4069_1;
wire na4070_1;
wire na4072_1;
wire na4072_4;
wire na4073_1;
wire na4073_4;
wire na4074_1;
wire na4075_1;
wire na4075_2;
wire na4075_4;
wire na4077_1;
wire na4078_1;
wire na4078_4;
wire na4079_1;
wire na4079_2;
wire na4079_4;
wire na4081_1;
wire na4081_2;
wire na4081_4;
wire na4083_1;
wire na4083_2;
wire na4085_1;
wire na4085_4;
wire na4087_1;
wire na4087_2;
wire na4087_4;
wire na4089_1;
wire na4089_2;
wire na4089_4;
wire na4091_1;
wire na4091_2;
wire na4091_4;
wire na4093_1;
wire na4093_2;
wire na4093_4;
wire na4095_1;
wire na4096_1;
wire na4096_2;
wire na4096_4;
wire na4098_1;
wire na4098_2;
wire na4098_4;
wire na4100_1;
wire na4100_2;
wire na4100_4;
wire na4102_1;
wire na4102_2;
wire na4102_4;
wire na4104_1;
wire na4104_2;
wire na4104_4;
wire na4105_1;
wire na4105_4;
wire na4106_1;
wire na4106_2;
wire na4106_4;
wire na4108_1;
wire na4108_2;
wire na4110_1;
wire na4110_4;
wire na4111_1;
wire na4111_2;
wire na4111_4;
wire na4113_1;
wire na4113_2;
wire na4116_1;
wire na4118_1;
wire na4118_1_i;
wire na4119_2;
wire na4119_2_i;
wire na4132_1;
wire na4132_1_i;
wire na4133_2;
wire na4133_2_i;
wire na4134_1;
wire na4134_1_i;
wire na4135_2;
wire na4135_2_i;
wire na4138_1;
wire na4138_1_i;
wire na4139_2;
wire na4139_2_i;
wire na4140_1;
wire na4140_1_i;
wire na4141_2;
wire na4141_2_i;
wire na4173_1;
wire na4173_1_i;
wire na4173_2;
wire na4173_2_i;
wire na4175_1;
wire na4175_1_i;
wire na4175_2;
wire na4175_2_i;
wire na4177_1;
wire na4177_1_i;
wire na4177_2;
wire na4177_2_i;
wire na4179_1;
wire na4179_1_i;
wire na4179_2;
wire na4179_2_i;
wire na4204_1;
wire na4204_1_i;
wire na4204_2;
wire na4204_2_i;
wire na4244_1;
wire na4244_1_i;
wire na4245_2;
wire na4245_2_i;
wire na4246_1;
wire na4246_1_i;
wire na4247_2;
wire na4247_2_i;
wire na4248_1;
wire na4248_1_i;
wire na4249_1;
wire na4249_1_i;
wire na4250_1;
wire na4250_1_i;
wire na4251_2;
wire na4251_2_i;
wire na4252_1;
wire na4252_1_i;
wire na4253_2;
wire na4253_2_i;
wire na4254_1;
wire na4254_1_i;
wire na4255_2;
wire na4255_2_i;
wire na4256_1;
wire na4256_1_i;
wire na4257_2;
wire na4257_2_i;
wire na4258_1;
wire na4258_1_i;
wire na4259_2;
wire na4259_2_i;
wire na4260_2;
wire na4260_2_i;
wire na4261_1;
wire na4261_1_i;
wire na4274_2;
wire na4274_2_i;
wire na4275_1;
wire na4275_1_i;
wire na4276_2;
wire na4276_2_i;
wire na4277_1;
wire na4277_1_i;
wire na4278_2;
wire na4278_2_i;
wire na4279_2;
wire na4279_2_i;
wire na4280_2;
wire na4280_2_i;
wire na4281_1;
wire na4281_1_i;
wire na4282_2;
wire na4282_2_i;
wire na4853_1;
wire na4853_1_i;
wire na4853_2;
wire na4853_2_i;
wire na4855_1;
wire na4855_1_i;
wire na4855_2;
wire na4855_2_i;
wire na4856_1;
wire na4856_1_i;
wire na4860_2;
wire na4860_2_i;
wire na4861_1;
wire na4861_1_i;
wire na4864_2;
wire na4864_2_i;
wire na4865_1;
wire na4865_1_i;
wire na4868_2;
wire na4868_2_i;
wire na4869_1;
wire na4869_1_i;
wire na4872_2;
wire na4872_2_i;
wire na4873_1;
wire na4873_1_i;
wire na4876_2;
wire na4876_2_i;
wire na4877_1;
wire na4877_1_i;
wire na4877_2;
wire na4877_2_i;
wire na4878_1;
wire na4878_1_i;
wire na4882_2;
wire na4882_2_i;
wire na4883_1;
wire na4883_1_i;
wire na4886_2;
wire na4886_2_i;
wire na4887_1;
wire na4887_1_i;
wire na4890_2;
wire na4890_2_i;
wire na4893_1;
wire na4893_1_i;
wire na4894_1;
wire na4894_1_i;
wire na4894_2;
wire na4894_2_i;
wire na4895_1;
wire na4895_1_i;
wire na4895_2;
wire na4895_2_i;
wire na4897_1;
wire na4897_1_i;
wire na4897_2;
wire na4897_2_i;
wire na4899_1;
wire na4899_1_i;
wire na4899_2;
wire na4899_2_i;
wire na4900_1;
wire na4900_1_i;
wire na4900_2;
wire na4900_2_i;
wire na4903_1;
wire na4903_1_i;
wire na4903_2;
wire na4903_2_i;
wire na4905_1;
wire na4905_1_i;
wire na4905_2;
wire na4905_2_i;
wire na4907_1;
wire na4907_1_i;
wire na4907_2;
wire na4907_2_i;
wire na4909_1;
wire na4909_1_i;
wire na4909_2;
wire na4909_2_i;
wire na4911_1;
wire na4911_1_i;
wire na4911_2;
wire na4911_2_i;
wire na4913_1;
wire na4913_1_i;
wire na4913_2;
wire na4913_2_i;
wire na4915_1;
wire na4915_1_i;
wire na4915_2;
wire na4915_2_i;
wire na4917_1;
wire na4917_1_i;
wire na4917_2;
wire na4917_2_i;
wire na4919_1;
wire na4919_1_i;
wire na4919_2;
wire na4919_2_i;
wire na4922_1;
wire na4922_1_i;
wire na4922_2;
wire na4922_2_i;
wire na4926_1;
wire na4926_1_i;
wire na4926_2;
wire na4926_2_i;
wire na4928_1;
wire na4928_1_i;
wire na4928_2;
wire na4928_2_i;
wire na4930_2;
wire na4930_2_i;
wire na4933_1;
wire na4933_1_i;
wire na4936_2;
wire na4936_2_i;
wire na5167_1;
wire na5167_1_i;
wire na5168_2;
wire na5168_2_i;
wire na5169_1;
wire na5169_1_i;
wire na5170_2;
wire na5170_2_i;
wire na5171_1;
wire na5171_1_i;
wire na5172_2;
wire na5172_2_i;
wire na5173_1;
wire na5173_1_i;
wire na5174_2;
wire na5174_2_i;
wire na5175_1;
wire na5175_1_i;
wire na5176_2;
wire na5176_2_i;
wire na5177_1;
wire na5177_1_i;
wire na5178_2;
wire na5178_2_i;
wire na5179_1;
wire na5179_1_i;
wire na5179_2;
wire na5179_2_i;
wire na5181_1;
wire na5181_1_i;
wire na5181_2;
wire na5181_2_i;
wire na5183_1;
wire na5183_1_i;
wire na5183_2;
wire na5183_2_i;
wire na5185_1;
wire na5185_1_i;
wire na5185_2;
wire na5185_2_i;
wire na5215_1;
wire na5215_1_i;
wire na5216_2;
wire na5216_2_i;
wire na5217_1;
wire na5217_1_i;
wire na5218_1;
wire na5218_1_i;
wire na5219_2;
wire na5219_2_i;
wire na5220_1;
wire na5220_1_i;
wire na5221_2;
wire na5221_2_i;
wire na5222_1;
wire na5222_1_i;
wire na5223_1;
wire na5223_1_i;
wire na5223_2;
wire na5223_2_i;
wire na5228_2;
wire na5228_2_i;
wire na5229_1;
wire na5229_1_i;
wire na5230_2;
wire na5230_2_i;
wire na5231_1;
wire na5231_1_i;
wire na5232_2;
wire na5232_2_i;
wire na5233_1;
wire na5233_1_i;
wire na5234_2;
wire na5234_2_i;
wire na5235_1;
wire na5235_1_i;
wire na5236_2;
wire na5236_2_i;
wire na5237_1;
wire na5237_1_i;
wire na5238_2;
wire na5238_2_i;
wire na5239_2;
wire na5239_2_i;
wire na5240_1;
wire na5240_1_i;
wire na5241_1;
wire na5241_1_i;
wire na5242_1;
wire na5242_1_i;
wire na5243_2;
wire na5243_2_i;
wire na5244_1;
wire na5244_1_i;
wire na5245_2;
wire na5245_2_i;
wire na5246_1;
wire na5246_1_i;
wire na5247_2;
wire na5247_2_i;
wire na5248_1;
wire na5248_1_i;
wire na5249_2;
wire na5249_2_i;
wire na5250_1;
wire na5250_1_i;
wire na5251_2;
wire na5251_2_i;
wire na5252_1;
wire na5252_1_i;
wire na5253_2;
wire na5253_2_i;
wire na5254_2;
wire na5254_2_i;
wire na5255_2;
wire na5255_2_i;
wire na5256_1;
wire na5256_1_i;
wire na5257_2;
wire na5257_2_i;
wire na5258_1;
wire na5258_1_i;
wire na5259_2;
wire na5259_2_i;
wire na5261_1;
wire na5261_1_i;
wire na5261_2;
wire na5261_2_i;
wire na5263_1;
wire na5263_1_i;
wire na5264_2;
wire na5264_2_i;
wire na5265_1;
wire na5265_1_i;
wire na5266_2;
wire na5266_2_i;
wire na5267_1;
wire na5267_1_i;
wire na5268_2;
wire na5268_2_i;
wire na5269_1;
wire na5269_1_i;
wire na5270_2;
wire na5270_2_i;
wire na5271_1;
wire na5271_1_i;
wire na5272_2;
wire na5272_2_i;
wire na5273_2;
wire na5273_2_i;
wire na5274_2;
wire na5274_2_i;
wire na5275_1;
wire na5275_1_i;
wire na5276_2;
wire na5276_2_i;
wire na5277_1;
wire na5277_1_i;
wire na5278_2;
wire na5278_2_i;
wire na5279_1;
wire na5279_1_i;
wire na5280_1;
wire na5280_1_i;
wire na5281_2;
wire na5281_2_i;
wire na5282_2;
wire na5282_2_i;
wire na5283_1;
wire na5283_1_i;
wire na5284_1;
wire na5284_1_i;
wire na5285_2;
wire na5285_2_i;
wire na5286_1;
wire na5286_1_i;
wire na5287_1;
wire na5287_1_i;
wire na5288_2;
wire na5288_2_i;
wire na5289_2;
wire na5289_2_i;
wire na5290_2;
wire na5290_2_i;
wire na5291_1;
wire na5291_1_i;
wire na5292_2;
wire na5292_2_i;
wire na5293_1;
wire na5293_1_i;
wire na5294_2;
wire na5294_2_i;
wire na5402_1;
wire na5402_1_i;
wire na5403_2;
wire na5403_2_i;
wire na5435_1;
wire na5435_1_i;
wire na5435_2;
wire na5435_2_i;
wire na5445_1;
wire na5445_1_i;
wire na5446_2;
wire na5446_2_i;
wire na5447_1;
wire na5447_1_i;
wire na5448_2;
wire na5448_2_i;
wire na5449_1;
wire na5449_1_i;
wire na5450_1;
wire na5450_1_i;
wire na5451_2;
wire na5451_2_i;
wire na5452_1;
wire na5452_1_i;
wire na5456_1;
wire na5456_1_i;
wire na5457_1;
wire na5457_1_i;
wire na5458_2;
wire na5458_2_i;
wire na5459_1;
wire na5459_1_i;
wire na5460_1;
wire na5460_1_i;
wire na5461_2;
wire na5461_2_i;
wire na5462_2;
wire na5462_2_i;
wire na5463_1;
wire na5463_1_i;
wire na5464_1;
wire na5464_1_i;
wire na5465_1;
wire na5465_1_i;
wire na5466_2;
wire na5466_2_i;
wire na5467_2;
wire na5467_2_i;
wire na5468_1;
wire na5468_1_i;
wire na5469_1;
wire na5469_1_i;
wire na5470_2;
wire na5470_2_i;
wire na5471_1;
wire na5471_1_i;
wire na5472_2;
wire na5472_2_i;
wire na5473_1;
wire na5473_1_i;
wire na5474_2;
wire na5474_2_i;
wire na5475_1;
wire na5475_1_i;
wire na5476_2;
wire na5476_2_i;
wire na5477_1;
wire na5477_1_i;
wire na5478_2;
wire na5478_2_i;
wire na5479_1;
wire na5479_1_i;
wire na5480_2;
wire na5480_2_i;
wire na5481_1;
wire na5481_1_i;
wire na5482_2;
wire na5482_2_i;
wire na5483_1;
wire na5483_1_i;
wire na5484_2;
wire na5484_2_i;
wire na5485_1;
wire na5485_1_i;
wire na5486_2;
wire na5486_2_i;
wire na5487_1;
wire na5487_1_i;
wire na5488_2;
wire na5488_2_i;
wire na5489_1;
wire na5489_1_i;
wire na5490_2;
wire na5490_2_i;
wire na5491_1;
wire na5491_1_i;
wire na5492_2;
wire na5492_2_i;
wire na5493_2;
wire na5493_2_i;
wire na5494_2;
wire na5494_2_i;
wire na5495_1;
wire na5495_1_i;
wire na5496_2;
wire na5496_2_i;
wire na5497_1;
wire na5497_1_i;
wire na5498_2;
wire na5498_2_i;
wire na5499_1;
wire na5499_1_i;
wire na5500_2;
wire na5500_2_i;
wire na5501_1;
wire na5501_1_i;
wire na5502_2;
wire na5502_2_i;
wire na5503_1;
wire na5503_1_i;
wire na5504_2;
wire na5504_2_i;
wire na5505_1;
wire na5505_1_i;
wire na5506_2;
wire na5506_2_i;
wire na5507_1;
wire na5507_1_i;
wire na5508_2;
wire na5508_2_i;
wire na5509_1;
wire na5509_1_i;
wire na5510_2;
wire na5510_2_i;
wire na5511_1;
wire na5511_1_i;
wire na5512_2;
wire na5512_2_i;
wire na5513_1;
wire na5513_1_i;
wire na5514_2;
wire na5514_2_i;
wire na5515_1;
wire na5515_1_i;
wire na5516_2;
wire na5516_2_i;
wire na5517_1;
wire na5517_1_i;
wire na5518_2;
wire na5518_2_i;
wire na5585_1;
wire na5585_1_i;
wire na5586_2;
wire na5586_2_i;
wire na5587_1;
wire na5587_1_i;
wire na5588_2;
wire na5588_2_i;
wire na5589_1;
wire na5589_1_i;
wire na5590_2;
wire na5590_2_i;
wire na5591_1;
wire na5591_1_i;
wire na5592_2;
wire na5592_2_i;
wire na5593_1;
wire na5593_1_i;
wire na5684_1;
wire na5684_1_i;
wire na5684_2;
wire na5684_2_i;
wire na5685_1;
wire na5685_1_i;
wire na5685_2;
wire na5685_2_i;
wire na5686_1;
wire na5686_1_i;
wire na5686_2;
wire na5686_2_i;
wire na5687_1;
wire na5687_1_i;
wire na5687_2;
wire na5687_2_i;
wire na5688_1;
wire na5688_1_i;
wire na5688_2;
wire na5688_2_i;
wire na5689_2;
wire na5689_2_i;
wire na5690_1;
wire na5690_1_i;
wire na5691_1;
wire na5691_1_i;
wire na5691_2;
wire na5691_2_i;
wire na5692_1;
wire na5692_1_i;
wire na5692_2;
wire na5692_2_i;
wire na5695_2;
wire na5695_2_i;
wire na5697_1;
wire na5697_1_i;
wire na5698_2;
wire na5698_2_i;
wire na5699_1;
wire na5699_1_i;
wire na5700_2;
wire na5700_2_i;
wire na5701_1;
wire na5701_1_i;
wire na5702_2;
wire na5702_2_i;
wire na5703_1;
wire na5703_1_i;
wire na5704_2;
wire na5704_2_i;
wire na5705_1;
wire na5705_1_i;
wire na5705_2;
wire na5705_2_i;
wire na5706_1;
wire na5706_1_i;
wire na5707_2;
wire na5707_2_i;
wire na5708_2;
wire na5708_2_i;
wire na5709_2;
wire na5709_2_i;
wire na5710_1;
wire na5710_1_i;
wire na5711_2;
wire na5711_2_i;
wire na5712_2;
wire na5712_2_i;
wire na5713_1;
wire na5713_1_i;
wire na5714_2;
wire na5714_2_i;
wire na5715_1;
wire na5715_1_i;
wire na5716_2;
wire na5716_2_i;
wire na5717_2;
wire na5717_2_i;
wire na5718_2;
wire na5718_2_i;
wire na5719_2;
wire na5719_2_i;
wire na5720_2;
wire na5720_2_i;
wire na5721_1;
wire na5721_1_i;
wire na5722_1;
wire na5722_1_i;
wire na5723_1;
wire na5723_1_i;
wire na5724_2;
wire na5724_2_i;
wire na5725_1;
wire na5725_1_i;
wire na5726_2;
wire na5726_2_i;
wire na5727_2;
wire na5727_2_i;
wire na5728_1;
wire na5728_1_i;
wire na5729_1;
wire na5729_1_i;
wire na5795_2;
wire na5795_2_i;
wire na5796_1;
wire na5796_1_i;
wire na5797_2;
wire na5797_2_i;
wire na5798_2;
wire na5798_2_i;
wire na5799_1;
wire na5799_1_i;
wire na5800_2;
wire na5800_2_i;
wire na5801_1;
wire na5801_1_i;
wire na5802_2;
wire na5802_2_i;
wire na5803_1;
wire na5803_1_i;
wire na5804_2;
wire na5804_2_i;
wire na5805_2;
wire na5805_2_i;
wire na5806_2;
wire na5806_2_i;
wire na5807_1;
wire na5807_1_i;
wire na5808_1;
wire na5808_1_i;
wire na5809_2;
wire na5809_2_i;
wire na5810_1;
wire na5810_1_i;
wire na5811_2;
wire na5811_2_i;
wire na5812_2;
wire na5812_2_i;
wire na5813_2;
wire na5813_2_i;
wire na5814_1;
wire na5814_1_i;
wire na5815_2;
wire na5815_2_i;
wire na5816_1;
wire na5816_1_i;
wire na5817_2;
wire na5817_2_i;
wire na5818_2;
wire na5818_2_i;
wire na5819_1;
wire na5819_1_i;
wire na5820_2;
wire na5820_2_i;
wire na5821_1;
wire na5821_1_i;
wire na5822_2;
wire na5822_2_i;
wire na5823_1;
wire na5823_1_i;
wire na5824_1;
wire na5824_1_i;
wire na5830_2;
wire na5830_2_i;
wire na5832_1;
wire na5832_1_i;
wire na5834_1;
wire na5834_1_i;
wire na5836_2;
wire na5836_2_i;
wire na5838_1;
wire na5838_1_i;
wire na5840_1;
wire na5840_1_i;
wire na5842_1;
wire na5842_1_i;
wire na5844_2;
wire na5844_2_i;
wire na5846_2;
wire na5846_2_i;
wire na5848_1;
wire na5848_1_i;
wire na5850_2;
wire na5850_2_i;
wire na5852_1;
wire na5852_1_i;
wire na5854_1;
wire na5854_1_i;
wire na5888_2;
wire na5888_2_i;
wire na5889_1;
wire na5889_1_i;
wire na5890_2;
wire na5890_2_i;
wire na5891_1;
wire na5891_1_i;
wire na5892_2;
wire na5892_2_i;
wire na5893_1;
wire na5893_1_i;
wire na5894_2;
wire na5894_2_i;
wire na5895_1;
wire na5895_1_i;
wire na5896_2;
wire na5896_2_i;
wire na5897_1;
wire na5897_1_i;
wire na5898_2;
wire na5898_2_i;
wire na5899_1;
wire na5899_1_i;
wire na5900_2;
wire na5900_2_i;
wire na5901_1;
wire na5901_1_i;
wire na5902_2;
wire na5902_2_i;
wire na5903_1;
wire na5903_1_i;
wire na5904_2;
wire na5904_2_i;
wire na5905_1;
wire na5905_1_i;
wire na5906_2;
wire na5906_2_i;
wire na5907_1;
wire na5907_1_i;
wire na5908_2;
wire na5908_2_i;
wire na5909_1;
wire na5909_1_i;
wire na5910_2;
wire na5910_2_i;
wire na5911_1;
wire na5911_1_i;
wire na5912_2;
wire na5912_2_i;
wire na5913_1;
wire na5913_1_i;
wire na5914_2;
wire na5914_2_i;
wire na5915_1;
wire na5915_1_i;
wire na5916_2;
wire na5916_2_i;
wire na5917_1;
wire na5917_1_i;
wire na5925_2;
wire na5925_2_i;
wire na5926_2;
wire na5926_2_i;
wire na5927_1;
wire na5927_1_i;
wire na5930_1;
wire na5930_1_i;
wire na5931_2;
wire na5931_2_i;
wire na5932_1;
wire na5932_1_i;
wire na5932_2;
wire na5932_2_i;
wire na5935_1;
wire na5935_1_i;
wire na5935_2;
wire na5935_2_i;
wire na5936_1;
wire na5936_1_i;
wire na5937_2;
wire na5937_2_i;
wire na5938_1;
wire na5938_1_i;
wire na5939_2;
wire na5939_2_i;
wire na5940_1;
wire na5940_1_i;
wire na5941_2;
wire na5941_2_i;
wire na5942_1;
wire na5942_1_i;
wire na5943_2;
wire na5943_2_i;
wire na5944_1;
wire na5944_1_i;
wire na5945_2;
wire na5945_2_i;
wire na5946_1;
wire na5946_1_i;
wire na5947_2;
wire na5947_2_i;
wire na5948_1;
wire na5948_1_i;
wire na5953_1;
wire na5953_1_i;
wire na5953_2;
wire na5953_2_i;
wire na5955_2;
wire na5955_2_i;
wire na5956_1;
wire na5956_1_i;
wire na5957_2;
wire na5957_2_i;
wire na5958_1;
wire na5958_1_i;
wire na5959_2;
wire na5959_2_i;
wire na5960_1;
wire na5960_1_i;
wire na5961_2;
wire na5961_2_i;
wire na5962_1;
wire na5962_1_i;
wire na5962_2;
wire na5962_2_i;
wire na5963_1;
wire na5963_1_i;
wire na5963_2;
wire na5963_2_i;
wire na5964_1;
wire na5964_1_i;
wire na5964_2;
wire na5964_2_i;
wire na5965_1;
wire na5965_1_i;
wire na5965_2;
wire na5965_2_i;
wire na5967_1;
wire na5967_1_i;
wire na5967_2;
wire na5967_2_i;
wire na5969_1;
wire na5969_1_i;
wire na5969_2;
wire na5969_2_i;
wire na5971_1;
wire na5971_1_i;
wire na5971_2;
wire na5971_2_i;
wire na5972_1;
wire na5972_1_i;
wire na5974_2;
wire na5974_2_i;
wire na5977_1;
wire na5977_1_i;
wire na5985_1;
wire na5985_1_i;
wire na6004_1;
wire na6004_1_i;
wire na6005_2;
wire na6005_2_i;
wire na6006_1;
wire na6006_1_i;
wire na6007_2;
wire na6007_2_i;
wire na6008_1;
wire na6008_1_i;
wire na6009_2;
wire na6009_2_i;
wire na6010_1;
wire na6010_1_i;
wire na6011_2;
wire na6011_2_i;
wire na6012_1;
wire na6012_1_i;
wire na6014_2;
wire na6014_2_i;
wire na6015_1;
wire na6015_1_i;
wire na6016_2;
wire na6016_2_i;
wire na6017_1;
wire na6017_1_i;
wire na6018_2;
wire na6018_2_i;
wire na6019_1;
wire na6019_1_i;
wire na6020_2;
wire na6020_2_i;
wire na6021_1;
wire na6021_1_i;
wire na6022_2;
wire na6022_2_i;
wire na6023_1;
wire na6023_1_i;
wire na6024_2;
wire na6024_2_i;
wire na6025_1;
wire na6025_1_i;
wire na6026_2;
wire na6026_2_i;
wire na6027_1;
wire na6027_1_i;
wire na6028_2;
wire na6028_2_i;
wire na6029_1;
wire na6029_1_i;
wire na6030_2;
wire na6030_2_i;
wire na6031_1;
wire na6031_1_i;
wire na6032_2;
wire na6032_2_i;
wire na6033_1;
wire na6033_1_i;
wire na6034_2;
wire na6034_2_i;
wire na6035_1;
wire na6035_1_i;
wire na6036_2;
wire na6036_2_i;
wire na6037_1;
wire na6037_1_i;
wire na6038_2;
wire na6038_2_i;
wire na6039_1;
wire na6039_1_i;
wire na6040_2;
wire na6040_2_i;
wire na6041_1;
wire na6041_1_i;
wire na6042_2;
wire na6042_2_i;
wire na6043_1;
wire na6043_1_i;
wire na6044_2;
wire na6044_2_i;
wire na6045_1;
wire na6045_1_i;
wire na6047_1;
wire na6047_1_i;
wire na6047_2;
wire na6047_2_i;
wire na6049_1;
wire na6049_1_i;
wire na6049_2;
wire na6049_2_i;
wire na6051_1;
wire na6051_1_i;
wire na6051_2;
wire na6051_2_i;
wire na6053_1;
wire na6053_1_i;
wire na6053_2;
wire na6053_2_i;
wire na6055_1;
wire na6055_1_i;
wire na6055_2;
wire na6055_2_i;
wire na6056_1;
wire na6056_4;
wire na6057_1;
wire na6057_1_i;
wire na6058_2;
wire na6058_2_i;
wire na6065_2;
wire na6065_2_i;
wire na6066_1;
wire na6066_1_i;
wire na6067_2;
wire na6067_2_i;
wire na6068_1;
wire na6068_1_i;
wire na6069_2;
wire na6069_2_i;
wire na6070_1;
wire na6070_1_i;
wire na6071_2;
wire na6071_2_i;
wire na6072_1;
wire na6072_1_i;
wire na6073_2;
wire na6073_2_i;
wire na6074_1;
wire na6074_1_i;
wire na6075_2;
wire na6075_2_i;
wire na6076_1;
wire na6076_1_i;
wire na6077_2;
wire na6077_2_i;
wire na6078_1;
wire na6078_1_i;
wire na6079_2;
wire na6079_2_i;
wire na6080_1;
wire na6080_1_i;
wire na6081_2;
wire na6081_2_i;
wire na6082_1;
wire na6082_1_i;
wire na6083_2;
wire na6083_2_i;
wire na6084_1;
wire na6084_1_i;
wire na6085_2;
wire na6085_2_i;
wire na6086_1;
wire na6086_1_i;
wire na6087_2;
wire na6087_2_i;
wire na6088_1;
wire na6088_1_i;
wire na6089_2;
wire na6089_2_i;
wire na6090_1;
wire na6090_1_i;
wire na6091_2;
wire na6091_2_i;
wire na6092_1;
wire na6092_1_i;
wire na6093_2;
wire na6093_2_i;
wire na6094_1;
wire na6094_1_i;
wire na6095_2;
wire na6095_2_i;
wire na6096_1;
wire na6096_1_i;
wire na6097_2;
wire na6097_2_i;
wire na6098_1;
wire na6098_1_i;
wire na6105_1;
wire na6105_1_i;
wire na6105_2;
wire na6105_2_i;
wire na6107_1;
wire na6107_1_i;
wire na6107_2;
wire na6107_2_i;
wire na6109_1;
wire na6109_1_i;
wire na6109_2;
wire na6109_2_i;
wire na6111_1;
wire na6111_1_i;
wire na6111_2;
wire na6111_2_i;
wire na6113_2;
wire na6113_2_i;
wire na6117_1;
wire na6117_1_i;
wire na6118_2;
wire na6118_2_i;
wire na6308_1;
wire na6308_1_i;
wire na6309_2;
wire na6309_2_i;
wire na6310_1;
wire na6310_1_i;
wire na6312_2;
wire na6312_2_i;
wire na6313_1;
wire na6313_1_i;
wire na6314_2;
wire na6314_2_i;
wire na6315_1;
wire na6315_1_i;
wire na6317_2;
wire na6317_2_i;
wire na6318_1;
wire na6318_1_i;
wire na6319_2;
wire na6319_2_i;
wire na6320_1;
wire na6320_1_i;
wire na6320_2;
wire na6320_2_i;
wire na6321_1;
wire na6321_1_i;
wire na6322_2;
wire na6322_2_i;
wire na6323_1;
wire na6323_1_i;
wire na6324_1;
wire na6324_1_i;
wire na6324_2;
wire na6324_2_i;
wire na6325_1;
wire na6325_1_i;
wire na6325_2;
wire na6325_2_i;
wire na6326_2;
wire na6326_2_i;
wire na6327_1;
wire na6327_1_i;
wire na6328_2;
wire na6328_2_i;
wire na6329_1;
wire na6329_1_i;
wire na6330_2;
wire na6330_2_i;
wire na6331_1;
wire na6331_1_i;
wire na6332_2;
wire na6332_2_i;
wire na6333_1;
wire na6333_1_i;
wire na6334_2;
wire na6334_2_i;
wire na6335_1;
wire na6335_1_i;
wire na6336_2;
wire na6336_2_i;
wire na6343_1;
wire na6343_4;
wire na6345_1;
wire na6345_2;
wire na6345_4;
wire na6347_1;
wire na6347_2;
wire na6347_4;
wire na6349_1;
wire na6349_2;
wire na6349_4;
wire na6351_1;
wire na6351_2;
wire na6351_4;
wire na6353_1;
wire na6353_2;
wire na6353_4;
wire na6354_1;
wire na6354_2;
wire na6354_4;
wire na6356_1;
wire na6356_2;
wire na6356_4;
wire na6358_1;
wire na6358_2;
wire na6358_4;
wire na6360_1;
wire na6360_2;
wire na6360_4;
wire na6362_1;
wire na6362_2;
wire na6362_4;
wire na6364_1;
wire na6364_2;
wire na6364_4;
wire na6367_1;
wire na6368_1;
wire na6368_2;
wire na6368_4;
wire na6370_1;
wire na6370_2;
wire na6370_4;
wire na6372_1;
wire na6372_2;
wire na6372_4;
wire na6374_1;
wire na6374_2;
wire na6374_4;
wire na6380_1;
wire na6380_4;
wire na6381_1;
wire na6381_2;
wire na6383_1;
wire na6384_1;
wire na6385_1;
wire na6386_1;
wire na6387_1;
wire na6388_1;
wire na6389_1;
wire na6390_1;
wire na6391_1;
wire na6392_1;
wire na6393_1;
wire na6394_1;
wire na6395_1;
wire na6396_1;
wire na6397_1;
wire na6398_1;
wire na6399_1;
wire na6400_1;
wire na6401_1;
wire na6402_1;
wire na6403_1;
wire na6404_1;
wire na6405_1;
wire na6406_1;
wire na6407_1;
wire na6408_1;
wire na6409_1;
wire na6410_1;
wire na6411_1;
wire na6412_1;
wire na6413_1;
wire na6414_1;
wire na6415_1;
wire na6416_1;
wire na6417_1;
wire na6418_1;
wire na6419_1;
wire na6420_1;
wire na6421_1;
wire na6422_1;
wire na6423_1;
wire na6424_1;
wire na6425_1;
wire na6426_1;
wire na6427_1;
wire na6428_1;
wire na6429_1;
wire na6430_1;
wire na6431_1;
wire na6432_1;
wire na6433_1;
wire na6434_1;
wire na6435_1;
wire na6436_1;
wire na6437_1;
wire na6438_1;
wire na6439_1;
wire na6440_1;
wire na6441_1;
wire na6442_1;
wire na6443_1;
wire na6444_1;
wire na6445_1;
wire na6446_1;
wire na6447_1;
wire na6447_1_i;
wire na6448_1;
wire na6448_1_i;
wire na6449_1;
wire na6449_1_i;
wire na6450_1;
wire na6450_1_i;
wire na6451_1;
wire na6451_1_i;
wire na6452_1;
wire na6452_1_i;
wire na6453_1;
wire na6453_1_i;
wire na6454_1;
wire na6455_1;
wire na6455_1_i;
wire na6456_1;
wire na6457_1;
wire na6457_1_i;
wire na6458_1;
wire na6458_1_i;
wire na6459_1;
wire na6460_1;
wire na6461_1;
wire na6461_1_i;
wire na6462_1;
wire na6462_1_i;
wire na6463_1;
wire na6464_1;
wire na6465_1;
wire na6465_1_i;
wire na6466_1;
wire na6467_1;
wire na6468_1;
wire na6469_1;
wire na6470_1;
wire na6471_1;
wire na6472_1;
wire na6473_1;
wire na6474_1;
wire na6475_1;
wire na6476_1;
wire na6477_1;
wire na6478_1;
wire na6479_1;
wire na6480_1;
wire na6481_1;
wire na6482_1;
wire na6483_1;
wire na6484_1;
wire na6485_1;
wire na6486_1;
wire na6487_1;
wire na6488_1;
wire na6489_1;
wire na6490_1;
wire na6491_1;
wire na6492_1;
wire na6493_1;
wire na6494_1;
wire na6495_1;
wire na6496_1;
wire na6497_1;
wire na6498_1;
wire na6498_1_i;
wire na6499_1;
wire na6499_1_i;
wire na6500_1;
wire na6500_1_i;
wire na6501_1;
wire na6501_1_i;
wire na6502_1;
wire na6502_1_i;
wire na6503_1;
wire na6503_1_i;
wire na6504_1;
wire na6504_1_i;
wire na6505_1;
wire na6505_1_i;
wire na6506_1;
wire na6506_1_i;
wire na6507_1;
wire na6507_1_i;
wire na6508_1;
wire na6508_1_i;
wire na6509_1;
wire na6509_1_i;
wire na6510_1;
wire na6510_1_i;
wire na6511_1;
wire na6511_1_i;
wire na6512_1;
wire na6512_1_i;
wire na6513_1;
wire na6513_1_i;
wire na6514_1;
wire na6514_1_i;
wire na6515_1;
wire na6515_1_i;
wire na6516_1;
wire na6516_1_i;
wire na6517_1;
wire na6517_1_i;
wire na6518_1;
wire na6518_1_i;
wire na6519_1;
wire na6519_1_i;
wire na6520_1;
wire na6520_1_i;
wire na6521_1;
wire na6521_1_i;
wire na6522_1;
wire na6522_1_i;
wire na6523_1;
wire na6523_1_i;
wire na6524_1;
wire na6524_1_i;
wire na6525_1;
wire na6525_1_i;
wire na6526_1;
wire na6526_1_i;
wire na6527_1;
wire na6527_1_i;
wire na6528_1;
wire na6528_1_i;
wire na6529_1;
wire na6529_1_i;
wire na6530_1;
wire na6531_1;
wire na6532_1;
wire na6533_1;
wire na6534_1;
wire na6535_1;
wire na6536_1;
wire na6537_1;
wire na6538_1;
wire na6539_1;
wire na6540_1;
wire na6541_1;
wire na6542_1;
wire na6543_1;
wire na6544_1;
wire na6545_1;
wire na6546_1;
wire na6547_1;
wire na6548_1;
wire na6549_1;
wire na6550_1;
wire na6551_1;
wire na6552_1;
wire na6553_1;
wire na6554_1;
wire na6555_1;
wire na6556_1;
wire na6557_1;
wire na6558_1;
wire na6559_1;
wire na6560_1;
wire na6561_1;
wire na6562_1;
wire na6562_4;
wire na6563_1;
wire na6563_2;
wire na6563_4;
wire na6565_1;
wire na6565_2;
wire na6565_4;
wire na6567_1;
wire na6567_2;
wire na6569_1;
wire na6570_1;
wire na6572_1;
wire na6573_1;
wire na6574_1;
wire na6575_1;
wire na6579_1;
wire na6580_1;
wire na6581_1;
wire na6582_1;
wire na6583_1;
wire na6584_1;
wire na6585_1;
wire na6586_1;
wire na6588_1;
wire na6590_1;
wire na6592_1;
wire na6593_1;
wire na6594_1;
wire na6595_1;
wire na6596_1;
wire na6597_1;
wire na6598_1;
wire na6599_1;
wire na6600_1;
wire na6601_1;
wire na6602_1;
wire na6604_1;
wire na6607_1;
wire na6611_1;
wire na6613_1;
wire na6615_1;
wire na6617_1;
wire na6624_1;
wire na6624_4;
wire na6626_1;
wire na6626_1_i;
wire na6626_2;
wire na6626_2_i;
wire na6627_2;
wire na6627_3;
wire na6627_4;
wire na6627_5;
wire na6627_6;
wire na6628_1;
wire na6630_1;
wire na6630_2;
wire na6630_3;
wire na6630_4;
wire na6630_5;
wire na6630_6;
wire na6630_7;
wire na6630_8;
wire na6630_9;
wire na6645_1;
wire na6645_2;
wire na6645_3;
wire na6645_4;
wire na6645_5;
wire na6645_6;
wire na6645_7;
wire na6645_8;
wire na6645_9;
wire na6646_2;
wire na6648_1;
wire na6648_2;
wire na6648_3;
wire na6648_4;
wire na6648_5;
wire na6648_6;
wire na6648_7;
wire na6648_8;
wire na6648_9;
wire na6649_2;
wire na6650_1;
wire na6650_2;
wire na6650_3;
wire na6650_4;
wire na6650_5;
wire na6650_6;
wire na6650_7;
wire na6650_8;
wire na6650_9;
wire na6651_1;
wire na6651_2;
wire na6651_3;
wire na6651_4;
wire na6651_5;
wire na6651_6;
wire na6651_7;
wire na6651_8;
wire na6651_9;
wire na6652_1;
wire na6652_9;
wire na6653_1;
wire na6653_2;
wire na6653_3;
wire na6653_4;
wire na6653_5;
wire na6653_6;
wire na6653_7;
wire na6653_8;
wire na6653_9;
wire na6654_2;
wire na6656_1;
wire na6656_9;
wire na6657_1;
wire na6657_2;
wire na6657_3;
wire na6657_4;
wire na6657_5;
wire na6657_6;
wire na6657_7;
wire na6657_8;
wire na6657_9;
wire na6658_2;
wire na6660_1;
wire na6660_9;
wire na6661_2;
wire na6662_1;
wire na6663_1;
wire na6664_1;
wire na6665_2;
wire na6666_2;
wire na6667_2;
wire na6668_1;
wire na6669_1;
wire na6669_9;
wire na6670_2;
wire na6671_2;
wire na6672_1;
wire na6673_1;
wire na6673_2;
wire na6674_2;
wire na6675_2;
wire na6676_1;
wire na6676_9;
wire na6677_2;
wire na6678_1;
wire na6679_2;
wire na6680_1;
wire na6680_9;
wire na6681_1;
wire na6682_2;
wire na6683_1;
wire na6683_9;
wire na6684_1;
wire na6684_2;
wire na6685_2;
wire na6686_1;
wire na6686_9;
wire na6687_2;
wire na6688_1;
wire na6688_9;
wire na6689_2;
wire na6690_1;
wire na6690_9;
wire na6691_2;
wire na6692_1;
wire na6693_1;
wire na6693_9;
wire na6694_2;
wire na6695_1;
wire na6696_1;
wire na6697_1;
wire na6697_9;
wire na6698_2;
wire na6699_2;
wire na6700_1;
wire na6700_2;
wire na6701_2;
wire na6702_1;
wire na6703_1;
wire na6703_9;
wire na6704_2;
wire na6705_1;
wire na6706_1;
wire na6707_1;
wire na6707_9;
wire na6708_2;
wire na6709_1;
wire na6710_1;
wire na6710_2;
wire na6711_1;
wire na6712_1;
wire na6713_1;
wire na6713_9;
wire na6714_2;
wire na6715_1;
wire na6715_9;
wire na6716_2;
wire na6716_2_i;
wire na6717_1;
wire na6717_1_i;
wire na6717_9;
wire na6718_2;
wire na6718_2_i;
wire na6719_1;
wire na6720_1;
wire na6720_1_i;
wire na6720_9;
wire na6721_2;
wire na6721_2_i;
wire na6722_1;
wire na6722_1_i;
wire na6722_9;
wire na6723_1;
wire na6724_1;
wire na6725_2;
wire na6725_2_i;
wire na6726_1;
wire na6726_1_i;
wire na6726_9;
wire na6727_1;
wire na6727_2;
wire na6728_2;
wire na6728_2_i;
wire na6729_1;
wire na6729_1_i;
wire na6729_9;
wire na6730_2;
wire na6730_2_i;
wire na6731_1;
wire na6731_1_i;
wire na6731_9;
wire na6732_2;
wire na6732_2_i;
wire na6733_1;
wire na6734_1;
wire na6734_1_i;
wire na6734_9;
wire na6735_2;
wire na6735_2_i;
wire na6736_2;
wire na6737_1;
wire na6737_1_i;
wire na6737_9;
wire na6738_2;
wire na6738_2_i;
wire na6739_1;
wire na6739_1_i;
wire na6739_9;
wire na6740_2;
wire na6740_2_i;
wire na6741_1;
wire na6742_1;
wire na6742_1_i;
wire na6742_9;
wire na6743_1;
wire na6744_2;
wire na6744_2_i;
wire na6745_1;
wire na6746_1;
wire na6746_1_i;
wire na6746_9;
wire na6747_2;
wire na6747_2_i;
wire na6748_1;
wire na6748_1_i;
wire na6748_9;
wire na6749_1;
wire na6750_1;
wire na6751_2;
wire na6751_2_i;
wire na6752_1;
wire na6753_1;
wire na6754_1;
wire na6754_1_i;
wire na6754_9;
wire na6755_2;
wire na6755_2_i;
wire na6756_1;
wire na6756_1_i;
wire na6756_9;
wire na6757_2;
wire na6757_2_i;
wire na6758_1;
wire na6758_1_i;
wire na6758_9;
wire na6759_1;
wire na6760_2;
wire na6760_2_i;
wire na6761_1;
wire na6761_1_i;
wire na6761_9;
wire na6762_2;
wire na6763_1;
wire na6763_9;
wire na6764_2;
wire na6765_1;
wire na6765_9;
wire na6766_2;
wire na6767_2;
wire na6768_1;
wire na6769_1;
wire na6770_1;
wire na6771_1;
wire na6772_1;
wire na6772_9;
wire na6773_2;
wire na6774_1;
wire na6775_1;
wire na6776_1;
wire na6777_2;
wire na6778_1;
wire na6778_2;
wire na6779_2;
wire na6780_2;
wire na6781_1;
wire na6782_2;
wire na6783_1;
wire na6784_1;
wire na6785_1;
wire na6785_9;
wire na6786_1;
wire na6787_1;
wire na6788_2;
wire na6789_1;
wire na6790_2;
wire na6791_2;
wire na6792_2;
wire na6793_2;
wire na6794_1;
wire na6795_1;
wire na6795_9;
wire na6796_2;
wire na6797_1;
wire na6798_2;
wire na6799_1;
wire na6800_2;
wire na6801_1;
wire na6801_9;
wire na6802_2;
wire na6803_1;
wire na6804_1;
wire na6804_9;
wire na6805_1;
wire na6806_2;
wire na6807_2;
wire na6808_1;
wire na6808_9;
wire na6809_2;
wire na6810_2;
wire na6811_1;
wire na6811_9;
wire na6812_1;
wire na6813_2;
wire na6814_1;
wire na6814_9;
wire na6815_2;
wire na6816_2;
wire na6817_1;
wire na6817_9;
wire na6818_2;
wire na6819_1;
wire na6819_9;
wire na6820_2;
wire na6821_1;
wire na6821_9;
wire na6822_2;
wire na6823_1;
wire na6824_1;
wire na6824_9;
wire na6825_2;
wire na6826_1;
wire na6826_9;
wire na6827_2;
wire na6828_1;
wire na6829_1;
wire na6829_9;
wire na6830_2;
wire na6831_1;
wire na6831_9;
wire na6832_2;
wire na6833_1;
wire na6833_9;
wire na6834_1;
wire na6835_2;
wire na6836_1;
wire na6837_1;
wire na6837_9;
wire na6838_2;
wire na6839_1;
wire na6839_2;
wire na6840_1;
wire na6840_9;
wire na6841_1;
wire na6842_2;
wire na6842_2_i;
wire na6843_1;
wire na6843_1_i;
wire na6843_9;
wire na6844_2;
wire na6844_2_i;
wire na6845_2;
wire na6846_1;
wire na6846_1_i;
wire na6846_9;
wire na6847_1;
wire na6848_2;
wire na6848_2_i;
wire na6849_1;
wire na6850_1;
wire na6850_1_i;
wire na6850_9;
wire na6851_2;
wire na6851_2_i;
wire na6852_1;
wire na6852_1_i;
wire na6852_9;
wire na6853_2;
wire na6854_2;
wire na6854_2_i;
wire na6855_1;
wire na6856_1;
wire na6856_1_i;
wire na6856_9;
wire na6857_2;
wire na6857_2_i;
wire na6858_1;
wire na6858_1_i;
wire na6858_9;
wire na6859_1;
wire na6860_2;
wire na6860_2_i;
wire na6861_1;
wire na6861_1_i;
wire na6861_9;
wire na6862_2;
wire na6862_2_i;
wire na6863_1;
wire na6863_1_i;
wire na6863_9;
wire na6864_1;
wire na6865_2;
wire na6865_2_i;
wire na6866_1;
wire na6867_1;
wire na6868_2;
wire na6869_2;
wire na6870_1;
wire na6871_1;
wire na6872_1;
wire na6872_1_i;
wire na6872_9;
wire na6873_2;
wire na6873_2_i;
wire na6874_1;
wire na6874_1_i;
wire na6874_9;
wire na6875_1;
wire na6876_2;
wire na6876_2_i;
wire na6877_1;
wire na6877_1_i;
wire na6877_9;
wire na6878_2;
wire na6878_2_i;
wire na6879_1;
wire na6880_1;
wire na6880_1_i;
wire na6880_9;
wire na6881_2;
wire na6882_2;
wire na6882_2_i;
wire na6883_1;
wire na6883_1_i;
wire na6883_9;
wire na6884_2;
wire na6884_2_i;
wire na6885_1;
wire na6885_1_i;
wire na6885_9;
wire na6886_1;
wire na6887_1;
wire na6888_1;
wire na6888_2;
wire na6889_2;
wire na6890_2;
wire na6890_2_i;
wire na6891_2;
wire na6892_1;
wire na6893_1;
wire na6893_1_i;
wire na6893_9;
wire na6894_2;
wire na6894_2_i;
wire na6895_1;
wire na6895_1_i;
wire na6895_9;
wire na6896_1;
wire na6897_2;
wire na6898_1;
wire na6898_9;
wire na6899_2;
wire na6900_1;
wire na6901_1;
wire na6901_9;
wire na6902_2;
wire na6903_1;
wire na6903_9;
wire na6904_1;
wire na6905_2;
wire na6906_1;
wire na6906_9;
wire na6907_1;
wire na6907_9;
wire na6908_2;
wire na6909_1;
wire na6910_1;
wire na6910_9;
wire na6911_2;
wire na6912_1;
wire na6912_9;
wire na6913_1;
wire na6914_2;
wire na6915_1;
wire na6915_9;
wire na6916_2;
wire na6917_1;
wire na6918_1;
wire na6918_9;
wire na6919_2;
wire na6920_1;
wire na6920_9;
wire na6921_1;
wire na6922_2;
wire na6923_1;
wire na6923_9;
wire na6924_2;
wire na6925_1;
wire na6926_1;
wire na6926_9;
wire na6927_2;
wire na6928_1;
wire na6928_9;
wire na6929_1;
wire na6930_2;
wire na6931_1;
wire na6931_9;
wire na6932_2;
wire na6933_1;
wire na6934_1;
wire na6934_9;
wire na6935_1;
wire na6936_1;
wire na6936_2;
wire na6937_2;
wire na6938_1;
wire na6939_2;
wire na6940_1;
wire na6940_9;
wire na6941_1;
wire na6942_1;
wire na6943_2;
wire na6944_1;
wire na6945_2;
wire na6946_1;
wire na6947_1;
wire na6948_1;
wire na6948_9;
wire na6949_2;
wire na6950_1;
wire na6951_1;
wire na6951_9;
wire na6952_2;
wire na6953_1;
wire na6953_9;
wire na6954_1;
wire na6955_2;
wire na6956_1;
wire na6956_9;
wire na6957_2;
wire na6958_1;
wire na6959_1;
wire na6959_9;
wire na6960_2;
wire na6961_1;
wire na6961_9;
wire na6962_1;
wire na6963_2;
wire na6964_1;
wire na6964_9;
wire na6965_2;
wire na6966_1;
wire na6967_1;
wire na6967_9;
wire na6968_2;
wire na6969_1;
wire na6969_9;
wire na6970_1;
wire na6971_2;
wire na6972_1;
wire na6972_9;
wire na6973_2;
wire na6974_1;
wire na6975_1;
wire na6975_9;
wire na6976_2;
wire na6977_1;
wire na6977_9;
wire na6978_1;
wire na6979_1;
wire na6980_1;
wire na6981_2;
wire na6982_1;
wire na6983_2;
wire na6984_1;
wire na6985_1;
wire na6985_9;
wire na6986_2;
wire na6987_1;
wire na6987_9;
wire na6988_1;
wire na6989_2;
wire na6990_1;
wire na6991_1;
wire na6991_9;
wire na6992_1;
wire na6993_2;
wire na6994_1;
wire na6994_9;
wire na6995_2;
wire na6996_1;
wire na6997_1;
wire na6998_1;
wire na6999_1;
wire na7000_2;
wire na7001_1;
wire na7002_1;
wire na7002_9;
wire na7003_1;
wire na7004_2;
wire na7005_2;
wire na7006_1;
wire na7007_1;
wire na7008_1;
wire na7009_1;
wire na7010_1;
wire na7011_1;
wire na7012_1;
wire na7012_9;
wire na7013_2;
wire na7014_1;
wire na7015_1;
wire na7016_1;
wire na7016_9;
wire na7017_1;
wire na7018_1;
wire na7019_1;
wire na7020_1;
wire na7021_1;
wire na7022_1;
wire na7023_1;
wire na7024_1;
wire na7025_1;
wire na7026_1;
wire na7027_1;
wire na7028_1;
wire na7029_1;
wire na7030_2;
wire na7031_1;
wire na7032_1;
wire na7033_2;
wire na7034_1;
wire na7035_1;
wire na7035_9;
wire na7036_1;
wire na7037_2;
wire na7038_2;
wire na7039_1;
wire na7040_2;
wire na7041_1;
wire na7042_2;
wire na7043_2;
wire na7044_2;
wire na7045_1;
wire na7045_9;
wire na7046_1;
wire na7047_1;
wire na7048_2;
wire na7049_2;
wire na7050_1;
wire na7050_9;
wire na7051_1;
wire na7052_2;
wire na7053_2;
wire na7054_1;
wire na7054_2;
wire na7055_1;
wire na7056_1;
wire na7056_9;
wire na7057_2;
wire na7058_2;
wire na7059_1;
wire na7060_1;
wire na7060_9;
wire na7061_1;
wire na7062_2;
wire na7063_1;
wire na7064_2;
wire na7065_1;
wire na7066_2;
wire na7067_1;
wire na7068_1;
wire na7069_1;
wire na7069_9;
wire na7070_2;
wire na7071_1;
wire na7072_1;
wire na7073_1;
wire na7073_9;
wire na7074_2;
wire na7075_1;
wire na7075_9;
wire na7076_1;
wire na7077_2;
wire na7078_1;
wire na7079_1;
wire na7079_9;
wire na7080_2;
wire na7081_1;
wire na7081_9;
wire na7082_1;
wire na7083_2;
wire na7084_1;
wire na7084_9;
wire na7085_2;
wire na7086_1;
wire na7087_1;
wire na7087_9;
wire na7088_2;
wire na7089_1;
wire na7089_9;
wire na7090_1;
wire na7091_2;
wire na7092_1;
wire na7092_9;
wire na7093_2;
wire na7094_1;
wire na7095_1;
wire na7095_9;
wire na7096_1;
wire na7097_1;
wire na7098_1;
wire na7099_2;
wire na7100_1;
wire na7101_1;
wire na7101_9;
wire na7102_2;
wire na7103_2;
wire na7104_1;
wire na7104_9;
wire na7105_1;
wire na7106_1;
wire na7107_2;
wire na7108_1;
wire na7109_1;
wire na7110_1;
wire na7111_1;
wire na7112_2;
wire na7113_1;
wire na7114_2;
wire na7115_1;
wire na7115_9;
wire na7116_2;
wire na7117_1;
wire na7117_9;
wire na7118_1;
wire na7119_2;
wire na7120_2;
wire na7121_1;
wire na7121_9;
wire na7122_1;
wire na7122_2;
wire na7123_2;
wire na7124_1;
wire na7125_1;
wire na7125_9;
wire na7126_2;
wire na7127_1;
wire na7127_9;
wire na7128_2;
wire na7129_1;
wire na7130_1;
wire na7130_9;
wire na7131_1;
wire na7132_2;
wire na7133_1;
wire na7134_1;
wire na7135_1;
wire na7136_1;
wire na7137_2;
wire na7138_1;
wire na7138_9;
wire na7139_2;
wire na7140_1;
wire na7141_1;
wire na7141_2;
wire na7142_2;
wire na7143_1;
wire na7143_9;
wire na7144_2;
wire na7145_1;
wire na7146_2;
wire na7147_1;
wire na7148_1;
wire na7149_2;
wire na7150_1;
wire na7150_9;
wire na7151_2;
wire na7152_1;
wire na7153_1;
wire na7153_9;
wire na7154_1;
wire na7155_2;
wire na7156_1;
wire na7156_9;
wire na7157_2;
wire na7158_1;
wire na7159_2;
wire na7160_1;
wire na7161_1;
wire na7162_1;
wire na7162_9;
wire na7163_2;
wire na7164_1;
wire na7165_1;
wire na7166_2;
wire na7167_1;
wire na7168_1;
wire na7168_9;
wire na7169_2;
wire na7170_1;
wire na7170_9;
wire na7171_1;
wire na7172_2;
wire na7173_1;
wire na7173_9;
wire na7174_2;
wire na7175_1;
wire na7175_9;
wire na7176_1;
wire na7177_2;
wire na7178_1;
wire na7179_1;
wire na7179_9;
wire na7180_2;
wire na7181_1;
wire na7181_9;
wire na7182_2;
wire na7183_1;
wire na7184_2;
wire na7185_1;
wire na7186_2;
wire na7187_1;
wire na7188_2;
wire na7189_1;
wire na7190_1;
wire na7191_1;
wire na7192_1;
wire na7193_2;
wire na7194_1;
wire na7194_9;
wire na7195_2;
wire na7196_1;
wire na7196_9;
wire na7197_2;
wire na7198_1;
wire na7199_1;
wire na7199_9;
wire na7200_2;
wire na7201_1;
wire na7201_9;
wire na7202_2;
wire na7203_1;
wire na7203_2;
wire na7204_1;
wire na7205_2;
wire na7206_2;
wire na7207_1;
wire na7208_1;
wire na7209_1;
wire na7210_1;
wire na7210_2;
wire na7211_1;
wire na7212_1;
wire na7213_1;
wire na7213_9;
wire na7214_2;
wire na7215_1;
wire na7215_9;
wire na7216_1;
wire na7217_1;
wire na7218_2;
wire na7219_1;
wire na7220_1;
wire na7221_2;
wire na7222_1;
wire na7223_1;
wire na7223_9;
wire na7224_1;
wire na7225_2;
wire na7226_1;
wire na7226_9;
wire na7227_2;
wire na7228_1;
wire na7229_1;
wire na7229_9;
wire na7230_2;
wire na7231_1;
wire na7231_9;
wire na7232_1;
wire na7233_1;
wire na7234_1;
wire na7235_1;
wire na7236_2;
wire na7237_1;
wire na7237_9;
wire na7238_2;
wire na7239_1;
wire na7239_9;
wire na7240_1;
wire na7241_2;
wire na7242_1;
wire na7242_9;
wire na7243_2;
wire na7244_1;
wire na7244_9;
wire na7245_1;
wire na7246_2;
wire na7247_1;
wire na7247_9;
wire na7248_2;
wire na7249_1;
wire na7249_9;
wire na7250_1;
wire na7251_2;
wire na7252_1;
wire na7252_9;
wire na7253_2;
wire na7254_1;
wire na7254_9;
wire na7255_1;
wire na7256_1;
wire na7257_2;
wire na7258_1;
wire na7259_2;
wire na7260_1;
wire na7261_1;
wire na7262_1;
wire na7262_2;
wire na7263_2;
wire na7264_1;
wire na7264_9;
wire na7265_1;
wire na7266_1;
wire na7267_2;
wire na7268_1;
wire na7268_9;
wire na7269_2;
wire na7270_1;
wire na7270_9;
wire na7271_1;
wire na7272_2;
wire na7273_1;
wire na7273_9;
wire na7274_2;
wire na7275_1;
wire na7275_9;
wire na7276_1;
wire na7277_2;
wire na7278_1;
wire na7278_2;
wire na7279_1;
wire na7280_2;
wire na7281_2;
wire na7282_1;
wire na7283_1;
wire na7283_9;
wire na7284_2;
wire na7285_1;
wire na7285_9;
wire na7286_1;
wire na7287_2;
wire na7288_1;
wire na7288_9;
wire na7289_2;
wire na7290_1;
wire na7291_2;
wire na7292_1;
wire na7293_1;
wire na7294_1;
wire na7295_2;
wire na7296_1;
wire na7297_2;
wire na7298_2;
wire na7299_2;
wire na7300_1;
wire na7301_1;
wire na7302_1;
wire na7302_9;
wire na7303_2;
wire na7304_1;
wire na7304_9;
wire na7305_1;
wire na7306_2;
wire na7307_1;
wire na7307_9;
wire na7308_2;
wire na7309_1;
wire na7309_9;
wire na7310_1;
wire na7311_1;
wire na7311_2;
wire na7312_2;
wire na7313_1;
wire na7314_1;
wire na7315_2;
wire na7316_1;
wire na7317_1;
wire na7318_2;
wire na7319_1;
wire na7320_2;
wire na7321_1;
wire na7322_1;
wire na7323_1;
wire na7324_2;
wire na7325_1;
wire na7326_1;
wire na7327_1;
wire na7328_2;
wire na7329_1;
wire na7330_1;
wire na7330_9;
wire na7331_2;
wire na7332_1;
wire na7332_9;
wire na7333_2;
wire na7334_1;
wire na7335_1;
wire na7336_1;
wire na7336_9;
wire na7337_2;
wire na7338_1;
wire na7338_9;
wire na7339_1;
wire na7340_2;
wire na7341_1;
wire na7341_9;
wire na7342_2;
wire na7343_2;
wire na7344_1;
wire na7344_2;
wire na7345_1;
wire na7345_2;
wire na7346_1;
wire na7347_1;
wire na7348_1;
wire na7349_1;
wire na7349_9;
wire na7350_2;
wire na7351_1;
wire na7351_9;
wire na7352_2;
wire na7353_1;
wire na7354_1;
wire na7355_1;
wire na7355_9;
wire na7356_2;
wire na7357_1;
wire na7357_9;
wire na7358_2;
wire na7359_1;
wire na7359_2;
wire na7360_1;
wire na7361_2;
wire na7362_2;
wire na7363_1;
wire na7364_1;
wire na7364_9;
wire na7365_2;
wire na7366_1;
wire na7366_9;
wire na7367_1;
wire na7368_2;
wire na7369_1;
wire na7369_9;
wire na7370_1;
wire na7371_1;
wire na7372_1;
wire na7373_2;
wire na7374_1;
wire na7375_2;
wire na7376_1;
wire na7377_1;
wire na7378_1;
wire na7378_9;
wire na7379_2;
wire na7380_1;
wire na7380_9;
wire na7381_1;
wire na7382_2;
wire na7383_1;
wire na7383_9;
wire na7384_2;
wire na7385_1;
wire na7386_1;
wire na7386_9;
wire na7387_2;
wire na7388_1;
wire na7388_9;
wire na7389_1;
wire na7390_2;
wire na7391_1;
wire na7391_9;
wire na7392_2;
wire na7393_1;
wire na7394_1;
wire na7394_9;
wire na7395_2;
wire na7396_1;
wire na7396_9;
wire na7397_1;
wire na7398_2;
wire na7399_1;
wire na7399_9;
wire na7400_2;
wire na7401_1;
wire na7402_1;
wire na7402_9;
wire na7403_2;
wire na7404_1;
wire na7404_9;
wire na7405_1;
wire na7406_2;
wire na7407_1;
wire na7407_9;
wire na7408_1;
wire na7409_1;
wire na7410_2;
wire na7411_1;
wire na7412_2;
wire na7413_1;
wire na7414_1;
wire na7415_1;
wire na7415_9;
wire na7416_2;
wire na7417_1;
wire na7418_1;
wire na7418_9;
wire na7419_2;
wire na7420_1;
wire na7420_9;
wire na7421_1;
wire na7422_2;
wire na7423_1;
wire na7423_9;
wire na7424_2;
wire na7425_1;
wire na7426_1;
wire na7426_9;
wire na7427_2;
wire na7428_1;
wire na7428_9;
wire na7429_1;
wire na7430_2;
wire na7431_1;
wire na7431_9;
wire na7432_2;
wire na7433_1;
wire na7434_1;
wire na7434_9;
wire na7435_2;
wire na7436_1;
wire na7436_9;
wire na7437_1;
wire na7438_2;
wire na7439_1;
wire na7439_9;
wire na7440_2;
wire na7441_1;
wire na7442_1;
wire na7442_9;
wire na7443_2;
wire na7444_1;
wire na7444_9;
wire na7445_1;
wire na7446_1;
wire na7447_2;
wire na7448_1;
wire na7449_1;
wire na7450_2;
wire na7451_1;
wire na7452_1;
wire na7452_9;
wire na7453_1;
wire na7454_2;
wire na7455_1;
wire na7455_9;
wire na7456_2;
wire na7457_1;
wire na7458_1;
wire na7458_9;
wire na7459_2;
wire na7460_1;
wire na7460_9;
wire na7461_1;
wire na7462_2;
wire na7463_1;
wire na7463_9;
wire na7464_2;
wire na7465_1;
wire na7466_1;
wire na7466_9;
wire na7467_2;
wire na7468_1;
wire na7468_9;
wire na7469_1;
wire na7470_2;
wire na7471_1;
wire na7471_9;
wire na7472_2;
wire na7473_1;
wire na7474_1;
wire na7474_9;
wire na7475_2;
wire na7476_1;
wire na7476_9;
wire na7477_1;
wire na7478_2;
wire na7479_1;
wire na7479_9;
wire na7480_2;
wire na7481_1;
wire na7482_1;
wire na7482_9;
wire na7483_1;
wire na7484_2;
wire na7485_1;
wire na7486_2;
wire na7487_2;
wire na7488_2;
wire na7489_1;
wire na7490_2;
wire na7491_1;
wire na7492_2;
wire na7493_1;
wire na7494_1;
wire na7495_2;
wire na7496_1;
wire na7497_1;
wire na7498_1;
wire na7498_9;
wire na7499_2;
wire na7500_1;
wire na7500_9;
wire na7501_1;
wire na7502_2;
wire na7503_1;
wire na7503_9;
wire na7504_2;
wire na7505_1;
wire na7506_1;
wire na7506_9;
wire na7507_2;
wire na7508_1;
wire na7508_9;
wire na7509_1;
wire na7510_2;
wire na7511_1;
wire na7511_9;
wire na7512_2;
wire na7513_1;
wire na7514_1;
wire na7514_9;
wire na7515_2;
wire na7516_1;
wire na7516_9;
wire na7517_1;
wire na7518_2;
wire na7519_1;
wire na7519_9;
wire na7520_2;
wire na7521_1;
wire na7522_1;
wire na7522_9;
wire na7523_2;
wire na7524_1;
wire na7524_9;
wire na7525_1;
wire na7526_2;
wire na7527_1;
wire na7527_9;
wire na7528_1;
wire na7529_1;
wire na7530_2;
wire na7531_1;
wire na7532_2;
wire na7533_1;
wire na7534_1;
wire na7535_1;
wire na7535_9;
wire na7536_2;
wire na7537_1;
wire na7538_2;
wire na7539_1;
wire na7539_9;
wire na7540_2;
wire na7541_1;
wire na7542_1;
wire na7542_9;
wire na7543_2;
wire na7544_1;
wire na7544_9;
wire na7545_1;
wire na7546_2;
wire na7547_1;
wire na7547_9;
wire na7548_2;
wire na7549_1;
wire na7550_1;
wire na7550_9;
wire na7551_2;
wire na7552_1;
wire na7552_9;
wire na7553_1;
wire na7554_2;
wire na7555_1;
wire na7555_9;
wire na7556_2;
wire na7557_1;
wire na7558_1;
wire na7558_9;
wire na7559_1;
wire na7559_9;
wire na7560_1;
wire na7560_9;
wire na7561_1;
wire na7562_2;
wire na7563_1;
wire na7563_9;
wire na7564_2;
wire na7565_1;
wire na7566_1;
wire na7566_9;
wire na7567_2;
wire na7567_2_i;
wire na7568_1;
wire na7568_1_i;
wire na7568_9;
wire na7569_1;
wire na7570_2;
wire na7570_2_i;
wire na7571_1;
wire na7571_1_i;
wire na7571_9;
wire na7572_2;
wire na7572_2_i;
wire na7573_1;
wire na7574_1;
wire na7574_1_i;
wire na7574_9;
wire na7575_2;
wire na7575_2_i;
wire na7576_1;
wire na7576_1_i;
wire na7576_9;
wire na7577_1;
wire na7578_2;
wire na7578_2_i;
wire na7579_1;
wire na7579_1_i;
wire na7579_9;
wire na7580_2;
wire na7580_2_i;
wire na7581_1;
wire na7582_1;
wire na7582_1_i;
wire na7582_9;
wire na7583_2;
wire na7583_2_i;
wire na7584_1;
wire na7584_1_i;
wire na7584_9;
wire na7585_1;
wire na7586_2;
wire na7586_2_i;
wire na7587_1;
wire na7587_1_i;
wire na7587_9;
wire na7588_2;
wire na7588_2_i;
wire na7589_1;
wire na7590_1;
wire na7590_1_i;
wire na7590_9;
wire na7591_2;
wire na7591_2_i;
wire na7592_1;
wire na7592_1_i;
wire na7592_9;
wire na7593_1;
wire na7594_2;
wire na7595_1;
wire na7596_1;
wire na7597_2;
wire na7598_1;
wire na7599_1;
wire na7600_2;
wire na7601_1;
wire na7602_2;
wire na7603_1;
wire na7603_9;
wire na7604_2;
wire na7605_1;
wire na7606_1;
wire na7606_9;
wire na7607_2;
wire na7608_1;
wire na7608_9;
wire na7609_1;
wire na7610_2;
wire na7611_1;
wire na7612_2;
wire na7613_2;
wire na7614_1;
wire na7615_1;
wire na7616_1;
wire na7617_1;
wire na7618_2;
wire na7619_1;
wire na7619_9;
wire na7620_2;
wire na7621_2;
wire na7622_1;
wire na7623_1;
wire na7624_1;
wire na7624_9;
wire na7625_2;
wire na7626_1;
wire na7626_9;
wire na7627_1;
wire na7628_2;
wire na7629_1;
wire na7629_2;
wire na7630_1;
wire na7631_2;
wire na7632_2;
wire na7633_1;
wire na7634_1;
wire na7634_9;
wire na7635_2;
wire na7636_1;
wire na7636_9;
wire na7637_1;
wire na7638_2;
wire na7639_1;
wire na7639_9;
wire na7640_2;
wire na7641_1;
wire na7642_1;
wire na7642_9;
wire na7643_1;
wire na7643_9;
wire na7644_1;
wire na7644_9;
wire na7645_1;
wire na7646_2;
wire na7647_2;
wire na7648_2;
wire na7649_1;
wire na7650_1;
wire na7650_9;
wire na7651_2;
wire na7652_1;
wire na7652_9;
wire na7653_1;
wire na7654_2;
wire na7655_1;
wire na7655_9;
wire na7656_2;
wire na7657_1;
wire na7658_1;
wire na7658_9;
wire na7659_2;
wire na7660_1;
wire na7660_9;
wire na7661_1;
wire na7662_2;
wire na7663_2;
wire na7664_2;
wire na7665_1;
wire na7666_2;
wire na7667_1;
wire na7668_2;
wire na7669_1;
wire na7670_2;
wire na7671_1;
wire na7672_1;
wire na7673_1;
wire na7674_2;
wire na7675_1;
wire na7676_2;
wire na7677_1;
wire na7678_2;
wire na7679_1;
wire na7680_2;
wire na7681_1;
wire na7682_2;
wire na7683_1;
wire na7684_2;
wire na7685_1;
wire na7686_2;
wire na7687_1;
wire na7688_1;
wire na7689_2;
wire na7690_2;
wire na7691_2;
wire na7692_1;
wire na7693_2;
wire na7694_1;
wire na7695_2;
wire na7696_1;
wire na7697_2;
wire na7698_1;
wire na7699_1;
wire na7700_1;
wire na7701_2;
wire na7702_1;
wire na7703_2;
wire na7704_1;
wire na7705_2;
wire na7706_1;
wire na7707_2;
wire na7708_2;
wire na7709_1;
wire na7710_2;
wire na7711_1;
wire na7711_9;
wire na7712_2;
wire na7713_1;
wire na7714_1;
wire na7714_9;
wire na7715_2;
wire na7716_1;
wire na7716_9;
wire na7717_2;
wire na7718_1;
wire na7718_9;
wire na7719_2;
wire na7720_1;
wire na7720_9;
wire na7721_2;
wire na7722_1;
wire na7722_9;
wire na7723_1;
wire na7724_2;
wire na7725_1;
wire na7725_9;
wire na7726_2;
wire na7727_1;
wire na7728_1;
wire na7729_2;
wire na7730_1;
wire na7731_1;
wire na7731_9;
wire na7732_1;
wire na7733_1;
wire na7734_2;
wire na7735_1;
wire na7736_1;
wire na7737_2;
wire na7738_1;
wire na7739_1;
wire na7739_9;
wire na7740_1;
wire na7741_1;
wire na7742_2;
wire na7743_2;
wire na7744_1;
wire na7744_9;
wire na7745_1;
wire na7746_1;
wire na7747_1;
wire na7748_1;
wire na7749_1;
wire na7750_2;
wire na7751_2;
wire na7752_1;
wire na7752_9;
wire na7753_1;
wire na7754_1;
wire na7755_1;
wire na7756_1;
wire na7757_1;
wire na7758_1;
wire na7758_9;
wire na7759_2;
wire na7760_1;
wire na7760_9;
wire na7761_1;
wire na7762_1;
wire na7763_1;
wire na7764_1;
wire na7765_1;
wire na7766_2;
wire na7767_2;
wire na7768_1;
wire na7768_9;
wire na7769_1;
wire na7770_1;
wire na7771_1;
wire na7772_1;
wire na7773_1;
wire na7774_1;
wire na7774_2;
wire na7775_1;
wire na7776_1;
wire na7777_2;
wire na7778_2;
wire na7779_1;
wire na7779_9;
wire na7780_1;
wire na7781_1;
wire na7782_1;
wire na7783_1;
wire na7783_9;
wire na7784_2;
wire na7785_1;
wire na7785_9;
wire na7786_1;
wire na7787_1;
wire na7788_1;
wire na7789_2;
wire na7790_1;
wire na7791_1;
wire na7791_9;
wire na7792_1;
wire na7793_1;
wire na7794_1;
wire na7795_2;
wire na7796_2;
wire na7797_1;
wire na7797_9;
wire na7798_1;
wire na7799_1;
wire na7800_1;
wire na7801_2;
wire na7801_2_i;
wire na7802_2;
wire na7803_1;
wire na7803_1_i;
wire na7803_9;
wire na7804_1;
wire na7805_1;
wire na7806_1;
wire na7807_2;
wire na7807_2_i;
wire na7808_2;
wire na7809_1;
wire na7809_1_i;
wire na7809_9;
wire na7810_1;
wire na7811_1;
wire na7812_1;
wire na7813_2;
wire na7813_2_i;
wire na7814_2;
wire na7815_1;
wire na7815_1_i;
wire na7815_9;
wire na7816_2;
wire na7817_1;
wire na7818_1;
wire na7819_2;
wire na7819_2_i;
wire na7820_2;
wire na7821_1;
wire na7821_1_i;
wire na7821_9;
wire na7822_1;
wire na7823_1;
wire na7824_1;
wire na7825_1;
wire na7826_2;
wire na7827_2;
wire na7827_2_i;
wire na7828_1;
wire na7829_1;
wire na7830_2;
wire na7831_1;
wire na7831_1_i;
wire na7831_9;
wire na7832_1;
wire na7833_1;
wire na7834_1;
wire na7835_2;
wire na7835_2_i;
wire na7836_1;
wire na7837_1;
wire na7838_2;
wire na7839_1;
wire na7839_1_i;
wire na7839_9;
wire na7840_1;
wire na7841_1;
wire na7842_1;
wire na7843_2;
wire na7843_2_i;
wire na7844_1;
wire na7845_1;
wire na7846_1;
wire na7847_1;
wire na7847_1_i;
wire na7847_9;
wire na7848_1;
wire na7849_1;
wire na7850_2;
wire na7851_2;
wire na7851_2_i;
wire na7852_1;
wire na7853_1;
wire na7854_1;
wire na7855_1;
wire na7855_1_i;
wire na7855_9;
wire na7856_1;
wire na7857_1;
wire na7858_2;
wire na7859_2;
wire na7859_2_i;
wire na7860_1;
wire na7861_1;
wire na7862_2;
wire na7863_1;
wire na7863_1_i;
wire na7863_9;
wire na7864_1;
wire na7865_1;
wire na7866_1;
wire na7867_2;
wire na7867_2_i;
wire na7868_1;
wire na7869_1;
wire na7870_2;
wire na7871_1;
wire na7871_1_i;
wire na7871_9;
wire na7872_1;
wire na7873_1;
wire na7874_2;
wire na7875_2;
wire na7875_2_i;
wire na7876_1;
wire na7877_1;
wire na7878_1;
wire na7879_1;
wire na7879_1_i;
wire na7879_9;
wire na7880_1;
wire na7881_1;
wire na7882_2;
wire na7883_2;
wire na7883_2_i;
wire na7884_1;
wire na7885_1;
wire na7886_1;
wire na7887_1;
wire na7887_1_i;
wire na7887_9;
wire na7888_1;
wire na7889_1;
wire na7890_2;
wire na7891_2;
wire na7892_2;
wire na7892_2_i;
wire na7893_1;
wire na7894_1;
wire na7894_1_i;
wire na7894_9;
wire na7895_1;
wire na7896_2;
wire na7896_2_i;
wire na7897_1;
wire na7898_1;
wire na7898_1_i;
wire na7898_9;
wire na7899_2;
wire na7900_2;
wire na7900_2_i;
wire na7901_1;
wire na7902_1;
wire na7902_1_i;
wire na7902_9;
wire na7903_1;
wire na7904_2;
wire na7904_2_i;
wire na7905_2;
wire na7906_1;
wire na7906_1_i;
wire na7906_9;
wire na7907_2;
wire na7907_2_i;
wire na7908_1;
wire na7908_1_i;
wire na7908_9;
wire na7909_2;
wire na7909_2_i;
wire na7910_1;
wire na7911_1;
wire na7911_1_i;
wire na7911_9;
wire na7912_1;
wire na7912_2;
wire na7913_2;
wire na7913_2_i;
wire na7914_1;
wire na7914_1_i;
wire na7914_9;
wire na7915_2;
wire na7915_2_i;
wire na7916_1;
wire na7916_1_i;
wire na7916_9;
wire na7917_2;
wire na7918_2;
wire na7919_1;
wire na7919_9;
wire na7920_2;
wire na7921_1;
wire na7921_9;
wire na7922_1;
wire na7923_2;
wire na7924_2;
wire na7925_1;
wire na7925_9;
wire na7926_1;
wire na7926_2;
wire na7927_2;
wire na7928_1;
wire na7929_1;
wire na7929_9;
wire na7930_2;
wire na7931_2;
wire na7932_1;
wire na7932_9;
wire na7933_2;
wire na7934_1;
wire na7934_2;
wire na7935_1;
wire na7935_9;
wire na7936_1;
wire na7937_2;
wire na7938_2;
wire na7939_1;
wire na7939_9;
wire na7940_2;
wire na7941_2;
wire na7942_2;
wire na7943_1;
wire na7943_9;
wire na7944_1;
wire na7945_2;
wire na7946_1;
wire na7946_9;
wire na7947_2;
wire na7948_1;
wire na7948_2;
wire na7949_1;
wire na7949_9;
wire na7950_2;
wire na7951_2;
wire na7952_2;
wire na7953_1;
wire na7953_2;
wire na7954_1;
wire na7955_1;
wire na7956_1;
wire na7956_9;
wire na7957_2;
wire na7958_2;
wire na7959_1;
wire na7960_1;
wire na7960_9;
wire na7961_1;
wire na7962_2;
wire na7963_1;
wire na7964_1;
wire na7964_9;
wire na7965_2;
wire na7966_1;
wire na7966_2;
wire na7967_1;
wire na7968_1;
wire na7968_9;
wire na7969_2;
wire na7970_1;
wire na7970_9;
wire na7971_1;
wire na7972_2;
wire na7973_1;
wire na7973_9;
wire na7974_2;
wire na7975_1;
wire na7976_1;
wire na7976_9;
wire na7977_2;
wire na7978_1;
wire na7978_9;
wire na7979_1;
wire na7980_2;
wire na7981_1;
wire na7981_9;
wire na7982_2;
wire na7983_1;
wire na7984_1;
wire na7984_9;
wire na7985_1;
wire na7985_9;
wire na7986_2;
wire na7987_1;
wire na7988_2;
wire na7989_1;
wire na7989_9;
wire na7990_2;
wire na7991_1;
wire na7991_9;
wire na7992_2;
wire na7993_1;
wire na7993_9;
wire na7994_2;
wire na7995_2;
wire na7996_1;
wire na7996_9;
wire na7997_1;
wire na7998_2;
wire na7999_1;
wire na7999_9;
wire na8000_1;
wire na8001_2;
wire na8002_1;
wire na8002_9;
wire na8003_1;
wire na8004_2;
wire na8005_1;
wire na8005_9;
wire na8006_2;
wire na8007_2;
wire na8008_1;
wire na8008_9;
wire na8009_1;
wire na8010_1;
wire na8010_9;
wire na8011_1;
wire na8011_9;
wire na8012_1;
wire na8013_2;
wire na8014_1;
wire na8014_9;
wire na8015_1;
wire na8016_2;
wire na8017_1;
wire na8017_9;
wire na8018_2;
wire na8019_2;
wire na8019_2_i;
wire na8020_1;
wire na8020_1_i;
wire na8020_9;
wire na8021_1;
wire na8022_2;
wire na8022_2_i;
wire na8023_1;
wire na8023_1_i;
wire na8023_9;
wire na8024_2;
wire na8025_2;
wire na8025_2_i;
wire na8026_1;
wire na8026_1_i;
wire na8026_9;
wire na8027_1;
wire na8028_2;
wire na8028_2_i;
wire na8029_1;
wire na8029_1_i;
wire na8029_9;
wire na8030_2;
wire na8031_2;
wire na8031_2_i;
wire na8032_1;
wire na8032_1_i;
wire na8032_9;
wire na8033_1;
wire na8034_2;
wire na8034_2_i;
wire na8035_1;
wire na8035_1_i;
wire na8035_9;
wire na8036_2;
wire na8037_2;
wire na8037_2_i;
wire na8038_1;
wire na8038_1_i;
wire na8038_9;
wire na8039_1;
wire na8040_2;
wire na8040_2_i;
wire na8041_1;
wire na8041_1_i;
wire na8041_9;
wire na8042_2;
wire na8042_2_i;
wire na8043_1;
wire na8043_1_i;
wire na8043_9;
wire na8044_2;
wire na8044_2_i;
wire na8045_1;
wire na8045_1_i;
wire na8045_9;
wire na8046_2;
wire na8047_1;
wire na8047_9;
wire na8048_2;
wire na8049_1;
wire na8049_9;
wire na8050_2;
wire na8051_1;
wire na8051_9;
wire na8052_2;
wire na8053_1;
wire na8053_9;
wire na8054_2;
wire na8055_1;
wire na8055_9;
wire na8056_2;
wire na8057_1;
wire na8057_9;
wire na8058_2;
wire na8059_2;
wire na8060_1;
wire na8060_9;
wire na8061_1;
wire na8062_2;
wire na8063_2;
wire na8064_1;
wire na8064_9;
wire na8065_2;
wire na8066_2;
wire na8067_2;
wire na8068_1;
wire na8068_9;
wire na8069_1;
wire na8070_2;
wire na8071_2;
wire na8072_1;
wire na8073_2;
wire na8074_1;
wire na8074_9;
wire na8075_2;
wire na8076_1;
wire na8077_2;
wire na8078_1;
wire na8079_1;
wire na8079_9;
wire na8080_1;
wire na8081_2;
wire na8082_1;
wire na8082_9;
wire na8083_2;
wire na8084_2;
wire na8085_1;
wire na8086_2;
wire na8087_1;
wire na8088_1;
wire na8088_9;
wire na8089_1;
wire na8090_2;
wire na8091_1;
wire na8092_2;
wire na8093_1;
wire na8094_1;
wire na8095_1;
wire na8096_2;
wire na8097_2;
wire na8098_1;
wire na8099_2;
wire na8100_1;
wire na8100_9;
wire na8101_1;
wire na8101_2;
wire na8102_2;
wire na8103_1;
wire na8104_1;
wire na8105_1;
wire na8105_9;
wire na8106_1;
wire na8107_1;
wire na8107_2;
wire na8108_2;
wire na8109_2;
wire na8110_1;
wire na8110_9;
wire na8111_2;
wire na8112_2;
wire na8113_1;
wire na8114_1;
wire na8114_9;
wire na8115_2;
wire na8116_2;
wire na8117_1;
wire na8117_9;
wire na8118_1;
wire na8119_2;
wire na8120_2;
wire na8121_1;
wire na8122_1;
wire na8122_9;
wire na8123_1;
wire na8124_2;
wire na8125_2;
wire na8126_1;
wire na8126_9;
wire na8127_2;
wire na8128_1;
wire na8128_9;
wire na8129_2;
wire na8130_1;
wire na8131_1;
wire na8131_9;
wire na8132_1;
wire na8132_2;
wire na8133_2;
wire na8134_2;
wire na8135_1;
wire na8135_9;
wire na8136_2;
wire na8137_1;
wire na8138_1;
wire na8138_9;
wire na8139_2;
wire na8140_1;
wire na8140_9;
wire na8141_2;
wire na8142_1;
wire na8143_1;
wire na8143_9;
wire na8144_2;
wire na8145_1;
wire na8145_9;
wire na8146_2;
wire na8147_1;
wire na8147_9;
wire na8148_1;
wire na8148_9;
wire na8149_1;
wire na8149_9;
wire na8150_2;
wire na8151_1;
wire na8152_2;
wire na8153_1;
wire na8153_9;
wire na8154_1;
wire na8155_2;
wire na8156_1;
wire na8156_9;
wire na8157_1;
wire na8157_9;
wire na8158_1;
wire na8159_1;
wire na8159_9;
wire na8160_2;
wire na8161_1;
wire na8161_9;
wire na8162_2;
wire na8163_1;
wire na8163_9;
wire na8164_2;
wire na8164_2_i;
wire na8165_1;
wire na8165_1_i;
wire na8165_9;
wire na8166_1;
wire na8167_2;
wire na8168_2;
wire na8168_2_i;
wire na8169_1;
wire na8169_1_i;
wire na8169_9;
wire na8170_2;
wire na8170_2_i;
wire na8171_1;
wire na8171_1_i;
wire na8171_9;
wire na8172_2;
wire na8172_2_i;
wire na8173_1;
wire na8174_2;
wire na8175_1;
wire na8176_1;
wire na8177_1;
wire na8178_1;
wire na8178_1_i;
wire na8178_9;
wire na8179_2;
wire na8179_2_i;
wire na8180_1;
wire na8180_1_i;
wire na8180_9;
wire na8181_2;
wire na8181_2_i;
wire na8182_1;
wire na8183_1;
wire na8184_2;
wire na8185_2;
wire na8186_1;
wire na8187_1;
wire na8188_1;
wire na8188_1_i;
wire na8188_9;
wire na8189_2;
wire na8189_2_i;
wire na8190_2;
wire na8191_1;
wire na8191_1_i;
wire na8191_9;
wire na8192_1;
wire na8192_2;
wire na8193_2;
wire na8193_2_i;
wire na8194_1;
wire na8194_1_i;
wire na8194_9;
wire na8195_2;
wire na8195_2_i;
wire na8196_1;
wire na8196_1_i;
wire na8196_9;
wire na8197_1;
wire na8198_2;
wire na8198_2_i;
wire na8199_1;
wire na8199_1_i;
wire na8199_9;
wire na8200_2;
wire na8200_2_i;
wire na8201_1;
wire na8201_1_i;
wire na8201_9;
wire na8202_2;
wire na8202_2_i;
wire na8203_1;
wire na8203_1_i;
wire na8203_9;
wire na8204_2;
wire na8204_2_i;
wire na8205_1;
wire na8205_1_i;
wire na8205_9;
wire na8206_2;
wire na8206_2_i;
wire na8207_1;
wire na8207_1_i;
wire na8207_9;
wire na8208_2;
wire na8208_2_i;
wire na8209_1;
wire na8209_1_i;
wire na8209_9;
wire na8210_2;
wire na8210_2_i;
wire na8211_1;
wire na8211_1_i;
wire na8211_9;
wire na8212_2;
wire na8212_2_i;
wire na8213_1;
wire na8213_1_i;
wire na8213_9;
wire na8214_2;
wire na8214_2_i;
wire na8215_1;
wire na8215_1_i;
wire na8215_9;
wire na8216_2;
wire na8216_2_i;
wire na8217_1;
wire na8217_1_i;
wire na8217_9;
wire na8218_2;
wire na8218_2_i;
wire na8219_1;
wire na8219_1_i;
wire na8219_9;
wire na8220_2;
wire na8221_1;
wire na8221_9;
wire na8222_2;
wire na8223_1;
wire na8223_9;
wire na8224_2;
wire na8225_1;
wire na8225_9;
wire na8226_2;
wire na8227_1;
wire na8227_9;
wire na8228_2;
wire na8229_1;
wire na8229_9;
wire na8230_2;
wire na8231_1;
wire na8231_9;
wire na8232_2;
wire na8233_1;
wire na8233_9;
wire na8234_2;
wire na8235_1;
wire na8235_9;
wire na8236_2;
wire na8237_1;
wire na8237_9;
wire na8238_2;
wire na8239_1;
wire na8239_9;
wire na8240_2;
wire na8241_1;
wire na8241_9;
wire na8242_2;
wire na8243_1;
wire na8243_9;
wire na8244_2;
wire na8245_1;
wire na8245_9;
wire na8246_2;
wire na8247_1;
wire na8247_9;
wire na8248_2;
wire na8249_1;
wire na8249_9;
wire na8250_2;
wire na8251_1;
wire na8251_9;
wire na8252_2;
wire na8253_1;
wire na8253_9;
wire na8254_2;
wire na8255_1;
wire na8255_9;
wire na8256_2;
wire na8257_1;
wire na8257_9;
wire na8258_2;
wire na8259_1;
wire na8259_9;
wire na8260_1;
wire na8260_9;
wire na8261_1;
wire na8261_9;
wire na8262_2;
wire na8263_2;
wire na8264_2;
wire na8265_1;
wire na8265_9;
wire na8266_2;
wire na8267_1;
wire na8268_1;
wire na8268_9;
wire na8269_2;
wire na8270_1;
wire na8270_9;
wire na8271_1;
wire na8272_1;
wire na8273_2;
wire na8274_2;
wire na8275_1;
wire na8275_2;
wire na8276_1;
wire na8276_9;
wire na8277_1;
wire na8277_2;
wire na8278_1;
wire na8278_2;
wire na8279_2;
wire na8280_1;
wire na8280_2;
wire na8281_1;
wire na8281_9;
wire na8282_2;
wire na8283_1;
wire na8283_2;
wire na8284_1;
wire na8284_9;
wire na8285_1;
wire na8285_2;
wire na8286_2;
wire na8287_1;
wire na8287_2;
wire na8288_1;
wire na8289_1;
wire na8289_2;
wire na8290_2;
wire na8291_1;
wire na8291_9;
wire na8292_1;
wire na8292_2;
wire na8293_2;
wire na8294_1;
wire na8294_2;
wire na8295_1;
wire na8295_2;
wire na8296_2;
wire na8297_1;
wire na8297_2;
wire na8298_1;
wire na8298_9;
wire na8299_2;
wire na8300_1;
wire na8301_1;
wire na8301_9;
wire na8302_1;
wire na8302_2;
wire na8303_2;
wire na8304_1;
wire na8304_2;
wire na8305_1;
wire na8306_1;
wire na8306_9;
wire na8307_1;
wire na8307_2;
wire na8308_2;
wire na8309_1;
wire na8309_2;
wire na8310_2;
wire na8311_1;
wire na8311_9;
wire na8312_1;
wire na8313_2;
wire na8314_1;
wire na8315_2;
wire na8316_2;
wire na8317_1;
wire na8318_1;
wire na8319_1;
wire na8320_1;
wire na8320_9;
wire na8321_2;
wire na8322_2;
wire na8323_1;
wire na8324_2;
wire na8325_2;
wire na8326_1;
wire na8326_9;
wire na8327_1;
wire na8328_2;
wire na8329_1;
wire na8330_1;
wire na8331_2;
wire na8332_2;
wire na8333_1;
wire na8334_1;
wire na8334_9;
wire na8335_2;
wire na8336_1;
wire na8336_9;
wire na8337_2;
wire na8338_1;
wire na8339_1;
wire na8340_2;
wire na8341_1;
wire na8342_1;
wire na8342_9;
wire na8343_1;
wire na8343_9;
wire na8344_1;
wire na8345_1;
wire na8346_1;
wire na8347_1;
wire na8347_9;
wire na8348_1;
wire na8349_2;
wire na8350_2;
wire na8351_1;
wire na8351_9;
wire na8352_1;
wire na8353_2;
wire na8354_1;
wire na8354_9;
wire na8355_2;
wire na8356_1;
wire na8356_9;
wire na8357_1;
wire na8357_2;
wire na8358_2;
wire na8359_1;
wire na8359_9;
wire na8360_1;
wire na8361_2;
wire na8362_2;
wire na8363_1;
wire na8364_2;
wire na8365_2;
wire na8366_1;
wire na8366_9;
wire na8367_1;
wire na8368_2;
wire na8369_1;
wire na8369_9;
wire na8370_1;
wire na8371_1;
wire na8371_2;
wire na8372_2;
wire na8373_1;
wire na8373_2;
wire na8374_2;
wire na8374_2_i;
wire na8375_1;
wire na8375_2;
wire na8376_1;
wire na8376_1_i;
wire na8376_9;
wire na8377_2;
wire na8378_1;
wire na8379_1;
wire na8380_2;
wire na8380_2_i;
wire na8381_1;
wire na8381_1_i;
wire na8381_9;
wire na8382_1;
wire na8383_2;
wire na8384_1;
wire na8384_2;
wire na8384_3;
wire na8384_3_i;
wire na8384_6;
wire na8385_1;
wire na8385_2;
wire na8385_3;
wire na8385_3_i;
wire na8385_6;
wire na8386_1;
wire na8386_2;
wire na8386_3;
wire na8386_3_i;
wire na8386_6;
wire na8387_1;
wire na8387_2;
wire na8387_3;
wire na8387_3_i;
wire na8387_6;
wire na8388_1;
wire na8388_2;
wire na8388_3;
wire na8388_3_i;
wire na8388_6;
wire na8389_1;
wire na8389_2;
wire na8389_3;
wire na8389_3_i;
wire na8389_6;
wire na8390_1;
wire na8390_2;
wire na8390_4;
wire na8390_7;
wire na8391_1;
wire na8391_3_i;
wire na8391_4;
wire na8391_5;
wire na8391_7;
wire na8392_3;
wire na8392_4;
wire na8392_5;
wire na8392_7;
wire na8393_1;
wire na8393_2;
wire na8393_3;
wire na8393_3_i;
wire na8393_4;
wire na8393_5;
wire na8393_7;
wire na8393_8;
wire na8394_1;
wire na8394_2;
wire na8394_4;
wire na8394_5;
wire na8394_7;
wire na8394_8;
wire na8395_3;
wire na8395_4;
wire na8395_5;
wire na8395_6;
wire na8395_7;
wire na8395_8;
wire na8396_3;
wire na8396_4;
wire na8396_5;
wire na8396_6;
wire na8396_7;
wire na8396_8;
wire na8397_3;
wire na8397_4;
wire na8397_5;
wire na8397_6;
wire na8397_7;
wire na8397_8;
wire na8398_3;
wire na8398_4;
wire na8398_5;
wire na8398_6;
wire na8398_7;
wire na8398_8;
wire na8399_3;
wire na8399_4;
wire na8399_5;
wire na8399_6;
wire na8399_7;
wire na8399_8;
wire na8400_2;
wire na8400_3;
wire na8400_3_i;
wire na8400_6;
wire na8401_1;
wire na8401_2;
wire na8401_4;
wire na8401_7;
wire na8402_1;
wire na8402_3_i;
wire na8402_4;
wire na8402_5;
wire na8402_7;
wire na8403_3;
wire na8403_4;
wire na8403_5;
wire na8403_7;
wire na8404_1;
wire na8404_2;
wire na8404_3;
wire na8404_3_i;
wire na8404_4;
wire na8404_5;
wire na8404_7;
wire na8404_8;
wire na8405_1;
wire na8405_2;
wire na8405_4;
wire na8405_5;
wire na8405_7;
wire na8405_8;
wire na8406_3;
wire na8406_4;
wire na8406_5;
wire na8406_6;
wire na8406_7;
wire na8406_8;
wire na8407_3;
wire na8407_4;
wire na8407_5;
wire na8407_6;
wire na8407_7;
wire na8407_8;
wire na8408_3;
wire na8408_4;
wire na8408_5;
wire na8408_6;
wire na8408_7;
wire na8408_8;
wire na8409_3;
wire na8409_4;
wire na8409_5;
wire na8409_6;
wire na8409_7;
wire na8409_8;
wire na8410_3;
wire na8410_4;
wire na8410_5;
wire na8410_6;
wire na8410_7;
wire na8410_8;
wire na8411_2;
wire na8411_3;
wire na8411_3_i;
wire na8411_6;
wire na8412_1;
wire na8412_2;
wire na8412_4;
wire na8412_7;
wire na8413_1;
wire na8413_3_i;
wire na8413_4;
wire na8413_5;
wire na8413_7;
wire na8414_4;
wire na8414_5;
wire na8414_7;
wire na8415_1;
wire na8415_2;
wire na8415_3_i;
wire na8415_4;
wire na8415_5;
wire na8415_7;
wire na8415_8;
wire na8416_1;
wire na8416_2;
wire na8416_4;
wire na8416_5;
wire na8416_7;
wire na8416_8;
wire na8417_1;
wire na8417_4;
wire na8417_5;
wire na8417_7;
wire na8417_8;
wire na8418_4;
wire na8418_5;
wire na8418_7;
wire na8418_8;
wire na8419_4;
wire na8419_5;
wire na8419_7;
wire na8419_8;
wire na8420_4;
wire na8420_5;
wire na8420_7;
wire na8420_8;
wire na8421_4;
wire na8421_5;
wire na8421_7;
wire na8421_8;
wire na8422_3_i;
wire na8423_2;
wire na8424_2;
wire na8425_2;
wire na8426_2;
wire na8427_2;
wire na8428_2;
wire na8429_2;
wire na8430_2;
wire na8431_2;
wire na8432_2;
wire na8433_2;
wire na8434_2;
wire na8435_2;
wire na8436_2;
wire na8437_2;
wire na8438_2;
wire na8439_2;
wire na8440_2;
wire na8441_2;
wire na8442_2;
wire na8443_2;
wire na8444_2;
wire na8445_2;
wire na8446_2;
wire na8447_2;
wire na8448_2;
wire na8449_2;
wire na8450_2;
wire na8451_2;
wire na8452_2;
wire na8453_2;
wire na8454_2;
wire na8455_2;
wire na8456_2;
wire na8457_2;
wire na8458_2;
wire na8459_2;
wire na8460_2;
wire na8461_2;
wire na8462_2;
wire na8463_2;
wire na8464_2;
wire na8465_2;
wire na8466_2;
wire na8467_2;
wire na8468_2;
wire na8469_2;
wire na8470_2;
wire na8471_2;
wire na8472_2;
wire na8473_2;
wire na8474_2;
wire na8475_2;
wire na8476_2;
wire na8477_2;
wire na8478_2;
wire na8479_2;
wire na8480_2;
wire na8481_2;
wire na8482_2;
wire na8483_2;
wire na8484_2;
wire na8485_2;
wire na8486_2;
wire na8487_2;
wire na8488_2;
wire na8489_2;
wire na8490_2;
wire na8491_2;
wire na8492_2;
wire na8493_2;
wire na8494_2;
wire na8495_2;
wire na8496_2;
wire na8497_2;
wire na8497_2_i;
wire na8498_1;
wire na8498_1_i;
wire na8498_9;
wire na8499_2;
wire na8499_2_i;
wire na8500_1;
wire na8500_1_i;
wire na8500_9;
wire na8501_2;
wire na8501_2_i;
wire na8502_1;
wire na8502_1_i;
wire na8502_9;
wire na8503_2;
wire na8503_2_i;
wire na8504_1;
wire na8504_1_i;
wire na8504_9;
wire na8505_2;
wire na8505_2_i;
wire na8506_1;
wire na8506_1_i;
wire na8506_9;
wire na8507_2;
wire na8507_2_i;
wire na8508_1;
wire na8508_1_i;
wire na8508_9;
wire na8509_2;
wire na8509_2_i;
wire na8510_1;
wire na8510_1_i;
wire na8510_9;
wire na8511_2;
wire na8511_2_i;
wire na8512_1;
wire na8512_1_i;
wire na8512_9;
wire na8513_2;
wire na8513_2_i;
wire na8514_1;
wire na8514_1_i;
wire na8514_9;
wire na8515_2;
wire na8515_2_i;
wire na8516_1;
wire na8516_1_i;
wire na8516_9;
wire na8517_2;
wire na8517_2_i;
wire na8518_1;
wire na8518_1_i;
wire na8518_9;
wire na8519_2;
wire na8519_2_i;
wire na8520_1;
wire na8520_1_i;
wire na8520_9;
wire na8521_2;
wire na8522_1;
wire na8522_9;
wire na8523_2;
wire na8524_1;
wire na8524_9;
wire na8525_2;
wire na8526_1;
wire na8526_9;
wire na8527_2;
wire na8528_1;
wire na8528_9;
wire na8529_2;
wire na8530_1;
wire na8530_9;
wire na8531_2;
wire na8532_1;
wire na8532_9;
wire na8533_2;
wire na8534_1;
wire na8534_9;
wire na8535_2;
wire na8536_1;
wire na8536_9;
wire na8537_2;
wire na8538_1;
wire na8538_9;
wire na8539_2;
wire na8540_1;
wire na8540_9;
wire na8541_1;
wire na8541_9;
wire na8542_1;
wire na8542_9;
wire na8543_2;
wire na8544_2;
wire na8545_2;
wire na8546_1;
wire na8546_9;
wire na8547_2;
wire na8548_1;
wire na8548_9;
wire na8549_2;
wire na8550_1;
wire na8550_9;
wire na8551_2;
wire na8552_1;
wire na8552_9;
wire na8553_2;
wire na8554_1;
wire na8554_9;
wire na8555_2;
wire na8556_1;
wire na8556_9;
wire na8557_2;
wire na8558_1;
wire na8558_9;
wire na8559_2;
wire na8560_1;
wire na8560_9;
wire na8561_2;
wire na8562_1;
wire na8562_9;
wire na8563_2;
wire na8564_1;
wire na8564_9;
wire na8565_2;
wire na8566_1;
wire na8566_9;
wire na8567_2;
wire na8568_1;
wire na8568_9;
wire na8569_2;
wire na8570_1;
wire na8570_9;
wire na8571_2;
wire na8572_1;
wire na8572_9;
wire na8573_2;
wire na8574_1;
wire na8574_9;
wire na8575_2;
wire na8576_1;
wire na8576_9;
wire na8577_1;
wire na8577_9;
wire na8578_1;
wire na8578_9;
wire na8579_2;
wire na8580_1;
wire na8580_9;
wire na8581_2;
wire na8582_1;
wire na8582_9;
wire na8583_1;
wire na8583_9;
wire na8584_1;
wire na8584_9;
wire na8585_2;
wire na8586_1;
wire na8586_9;
wire na8587_2;
wire na8588_1;
wire na8588_9;
wire na8589_2;
wire na8589_2_i;
wire na8590_1;
wire na8590_1_i;
wire na8590_9;
wire na8591_2;
wire na8591_2_i;
wire na8592_1;
wire na8592_1_i;
wire na8592_9;
wire na8593_2;
wire na8593_2_i;
wire na8594_1;
wire na8594_1_i;
wire na8594_9;
wire na8595_2;
wire na8595_2_i;
wire na8596_1;
wire na8596_1_i;
wire na8596_9;
wire na8597_2;
wire na8597_2_i;
wire na8598_1;
wire na8598_1_i;
wire na8598_9;
wire na8599_2;
wire na8599_2_i;
wire na8600_1;
wire na8600_1_i;
wire na8600_9;
wire na8601_2;
wire na8601_2_i;
wire na8602_1;
wire na8602_1_i;
wire na8602_9;
wire na8603_2;
wire na8603_2_i;
wire na8604_1;
wire na8604_1_i;
wire na8604_9;
wire na8605_2;
wire na8605_2_i;
wire na8606_1;
wire na8606_1_i;
wire na8606_9;
wire na8607_2;
wire na8607_2_i;
wire na8608_1;
wire na8608_1_i;
wire na8608_9;
wire na8609_2;
wire na8609_2_i;
wire na8610_1;
wire na8610_1_i;
wire na8610_9;
wire na8611_2;
wire na8611_2_i;
wire na8612_1;
wire na8612_1_i;
wire na8612_9;
wire na8613_2;
wire na8613_2_i;
wire na8614_1;
wire na8614_1_i;
wire na8614_9;
wire na8615_2;
wire na8615_2_i;
wire na8616_1;
wire na8616_1_i;
wire na8616_9;
wire na8617_2;
wire na8617_2_i;
wire na8618_1;
wire na8618_1_i;
wire na8618_9;
wire na8619_2;
wire na8619_2_i;
wire na8620_1;
wire na8620_1_i;
wire na8620_9;
wire na8621_2;
wire na8621_2_i;
wire na8622_1;
wire na8622_1_i;
wire na8622_9;
wire na8623_2;
wire na8623_2_i;
wire na8624_1;
wire na8624_1_i;
wire na8624_9;
wire na8625_2;
wire na8625_2_i;
wire na8626_1;
wire na8626_1_i;
wire na8626_9;
wire na8627_2;
wire na8627_2_i;
wire na8628_1;
wire na8628_1_i;
wire na8628_9;
wire na8629_2;
wire na8630_1;
wire na8630_9;
wire na8631_2;
wire na8632_1;
wire na8632_9;
wire na8633_2;
wire na8634_1;
wire na8634_9;
wire na8635_2;
wire na8636_1;
wire na8636_9;
wire na8637_2;
wire na8638_1;
wire na8638_9;
wire na8639_2;
wire na8640_1;
wire na8640_9;
wire na8641_2;
wire na8642_1;
wire na8642_9;
wire na8643_2;
wire na8644_1;
wire na8644_9;
wire na8645_2;
wire na8646_1;
wire na8646_9;
wire na8647_2;
wire na8648_1;
wire na8648_9;
wire na8649_2;
wire na8650_1;
wire na8650_9;
wire na8651_2;
wire na8652_1;
wire na8652_9;
wire na8653_2;
wire na8654_1;
wire na8654_9;
wire na8655_2;
wire na8656_1;
wire na8656_9;
wire na8657_2;
wire na8658_1;
wire na8658_9;
wire na8659_2;
wire na8660_1;
wire na8660_9;
wire na8661_2;
wire na8662_1;
wire na8662_9;
wire na8663_2;
wire na8664_1;
wire na8664_9;
wire na8665_2;
wire na8666_1;
wire na8666_9;
wire na8667_2;
wire na8668_1;
wire na8668_9;
wire na8669_1;
wire na8669_9;
wire na8670_1;
wire na8670_9;
wire na8671_2;
wire na8672_2;
wire na8673_2;
wire na8674_1;
wire na8674_9;
wire na8675_2;
wire na8676_1;
wire na8676_9;
wire na8677_2;
wire na8678_1;
wire na8678_9;
wire na8679_2;
wire na8680_1;
wire na8680_9;
wire na8681_2;
wire na8682_1;
wire na8682_9;
wire na8683_2;
wire na8684_1;
wire na8684_9;
wire na8685_2;
wire na8686_1;
wire na8686_9;
wire na8687_2;
wire na8688_1;
wire na8688_9;
wire na8689_2;
wire na8690_1;
wire na8690_9;
wire na8691_2;
wire na8692_1;
wire na8692_9;
wire na8693_2;
wire na8694_1;
wire na8694_9;
wire na8695_2;
wire na8696_1;
wire na8696_9;
wire na8697_2;
wire na8698_1;
wire na8698_9;
wire na8699_2;
wire na8700_1;
wire na8700_9;
wire na8701_2;
wire na8702_1;
wire na8702_9;
wire na8703_2;
wire na8704_1;
wire na8704_9;
wire na8705_1;
wire na8705_9;
wire na8706_1;
wire na8706_9;
wire na8707_2;
wire na8708_1;
wire na8708_9;
wire na8709_2;
wire na8710_1;
wire na8710_9;
wire na8711_1;
wire na8711_9;
wire na8712_1;
wire na8712_9;
wire na8713_2;
wire na8714_1;
wire na8714_9;
wire na8715_2;
wire na8716_1;
wire na8716_9;
wire na8717_2;
wire na8717_2_i;
wire na8718_1;
wire na8718_1_i;
wire na8718_9;
wire na8719_2;
wire na8719_2_i;
wire na8720_1;
wire na8720_1_i;
wire na8720_9;
wire na8721_2;
wire na8721_2_i;
wire na8722_1;
wire na8722_1_i;
wire na8722_9;
wire na8723_2;
wire na8723_2_i;
wire na8724_1;
wire na8724_1_i;
wire na8724_9;
wire na8725_2;
wire na8725_2_i;
wire na8726_1;
wire na8726_1_i;
wire na8726_9;
wire na8727_2;
wire na8727_2_i;
wire na8728_1;
wire na8728_1_i;
wire na8728_9;
wire na8729_2;
wire na8729_2_i;
wire na8730_1;
wire na8730_1_i;
wire na8730_9;
wire na8731_2;
wire na8731_2_i;
wire na8732_1;
wire na8732_1_i;
wire na8732_9;
wire na8733_2;
wire na8733_2_i;
wire na8734_1;
wire na8734_1_i;
wire na8734_9;
wire na8735_2;
wire na8735_2_i;
wire na8736_1;
wire na8736_1_i;
wire na8736_9;
wire na8737_2;
wire na8737_2_i;
wire na8738_1;
wire na8738_1_i;
wire na8738_9;
wire na8739_2;
wire na8739_2_i;
wire na8740_1;
wire na8740_1_i;
wire na8740_9;
wire na8741_2;
wire na8741_2_i;
wire na8742_1;
wire na8742_1_i;
wire na8742_9;
wire na8743_2;
wire na8743_2_i;
wire na8744_1;
wire na8744_1_i;
wire na8744_9;
wire na8745_2;
wire na8745_2_i;
wire na8746_1;
wire na8746_1_i;
wire na8746_9;
wire na8747_2;
wire na8747_2_i;
wire na8748_1;
wire na8748_1_i;
wire na8748_9;
wire na8749_2;
wire na8749_2_i;
wire na8750_1;
wire na8750_1_i;
wire na8750_9;
wire na8751_2;
wire na8751_2_i;
wire na8752_1;
wire na8752_1_i;
wire na8752_9;
wire na8753_2;
wire na8753_2_i;
wire na8754_1;
wire na8754_1_i;
wire na8754_9;
wire na8755_2;
wire na8755_2_i;
wire na8756_1;
wire na8756_1_i;
wire na8756_9;
wire na8757_2;
wire na8758_1;
wire na8758_9;
wire na8759_2;
wire na8760_1;
wire na8760_9;
wire na8761_2;
wire na8762_1;
wire na8762_9;
wire na8763_2;
wire na8764_1;
wire na8764_9;
wire na8765_2;
wire na8766_1;
wire na8766_9;
wire na8767_2;
wire na8768_1;
wire na8768_9;
wire na8769_2;
wire na8770_1;
wire na8770_9;
wire na8771_2;
wire na8772_1;
wire na8772_9;
wire na8773_2;
wire na8774_1;
wire na8774_9;
wire na8775_2;
wire na8776_1;
wire na8776_9;
wire na8777_2;
wire na8778_1;
wire na8778_9;
wire na8779_2;
wire na8780_1;
wire na8780_9;
wire na8781_2;
wire na8782_1;
wire na8782_9;
wire na8783_2;
wire na8784_1;
wire na8784_9;
wire na8785_2;
wire na8786_1;
wire na8786_9;
wire na8787_2;
wire na8788_1;
wire na8788_9;
wire na8789_2;
wire na8790_1;
wire na8790_9;
wire na8791_2;
wire na8792_1;
wire na8792_9;
wire na8793_2;
wire na8794_1;
wire na8794_9;
wire na8795_2;
wire na8796_1;
wire na8796_9;
wire na8797_1;
wire na8797_9;
wire na8798_2;
wire na8799_2;
wire na8800_1;
wire na8800_9;
wire na8801_2;
wire na8802_1;
wire na8802_9;
wire na8803_2;
wire na8804_1;
wire na8804_9;
wire na8805_2;
wire na8806_1;
wire na8806_9;
wire na8807_2;
wire na8808_1;
wire na8808_9;
wire na8809_2;
wire na8810_1;
wire na8810_9;
wire na8811_2;
wire na8812_1;
wire na8812_9;
wire na8813_2;
wire na8814_1;
wire na8814_9;
wire na8815_1;
wire na8815_9;
wire na8816_1;
wire na8816_9;
wire na8817_2;
wire na8818_1;
wire na8818_9;
wire na8819_2;
wire na8820_1;
wire na8820_9;
wire na8821_2;
wire na8821_2_i;
wire na8822_1;
wire na8822_1_i;
wire na8822_9;
wire na8823_2;
wire na8823_2_i;
wire na8824_1;
wire na8824_1_i;
wire na8824_9;
wire na8825_2;
wire na8825_2_i;
wire na8826_1;
wire na8826_1_i;
wire na8826_9;
wire na8827_2;
wire na8827_2_i;
wire na8828_1;
wire na8828_1_i;
wire na8828_9;
wire na8829_2;
wire na8829_2_i;
wire na8830_1;
wire na8830_1_i;
wire na8830_9;
wire na8831_2;
wire na8831_2_i;
wire na8832_1;
wire na8832_1_i;
wire na8832_9;
wire na8833_2;
wire na8833_2_i;
wire na8834_1;
wire na8834_1_i;
wire na8834_9;
wire na8835_2;
wire na8835_2_i;
wire na8836_1;
wire na8836_1_i;
wire na8836_9;
wire na8837_2;
wire na8837_2_i;
wire na8838_1;
wire na8838_1_i;
wire na8838_9;
wire na8839_2;
wire na8839_2_i;
wire na8840_1;
wire na8840_1_i;
wire na8840_9;
wire na8841_2;
wire na8842_1;
wire na8842_9;
wire na8843_2;
wire na8844_1;
wire na8844_9;
wire na8845_2;
wire na8846_1;
wire na8846_9;
wire na8847_2;
wire na8848_1;
wire na8848_9;
wire na8849_2;
wire na8850_1;
wire na8850_9;
wire na8851_2;
wire na8852_1;
wire na8852_9;
wire na8853_2;
wire na8854_1;
wire na8854_9;
wire na8855_2;
wire na8856_1;
wire na8856_9;
wire na8857_2;
wire na8858_1;
wire na8858_9;
wire na8859_2;
wire na8860_1;
wire na8860_9;
wire na8861_1;
wire na8861_9;
wire na8862_1;
wire na8862_9;
wire na8863_2;
wire na8864_2;
wire na8865_2;
wire na8866_1;
wire na8866_9;
wire na8867_2;
wire na8868_1;
wire na8868_9;
wire na8869_2;
wire na8870_1;
wire na8870_9;
wire na8871_2;
wire na8872_1;
wire na8872_9;
wire na8873_2;
wire na8874_1;
wire na8874_9;
wire na8875_2;
wire na8876_1;
wire na8876_9;
wire na8877_2;
wire na8878_1;
wire na8878_9;
wire na8879_2;
wire na8880_1;
wire na8880_9;
wire na8881_2;
wire na8882_1;
wire na8882_9;
wire na8883_2;
wire na8884_1;
wire na8884_9;
wire na8885_2;
wire na8886_1;
wire na8886_9;
wire na8887_2;
wire na8888_1;
wire na8888_9;
wire na8889_2;
wire na8890_1;
wire na8890_9;
wire na8891_2;
wire na8892_1;
wire na8892_9;
wire na8893_2;
wire na8894_1;
wire na8894_9;
wire na8895_2;
wire na8896_1;
wire na8896_9;
wire na8897_1;
wire na8897_9;
wire na8898_1;
wire na8898_9;
wire na8899_2;
wire na8900_1;
wire na8900_9;
wire na8901_2;
wire na8902_1;
wire na8902_9;
wire na8903_1;
wire na8903_9;
wire na8904_1;
wire na8904_9;
wire na8905_2;
wire na8906_1;
wire na8906_9;
wire na8907_2;
wire na8908_1;
wire na8908_9;
wire na8909_2;
wire na8909_2_i;
wire na8910_1;
wire na8910_1_i;
wire na8910_9;
wire na8911_2;
wire na8911_2_i;
wire na8912_1;
wire na8912_1_i;
wire na8912_9;
wire na8913_2;
wire na8913_2_i;
wire na8914_1;
wire na8914_1_i;
wire na8914_9;
wire na8915_2;
wire na8915_2_i;
wire na8916_1;
wire na8916_1_i;
wire na8916_9;
wire na8917_2;
wire na8917_2_i;
wire na8918_1;
wire na8918_1_i;
wire na8918_9;
wire na8919_2;
wire na8919_2_i;
wire na8920_1;
wire na8920_1_i;
wire na8920_9;
wire na8921_2;
wire na8921_2_i;
wire na8922_1;
wire na8922_1_i;
wire na8922_9;
wire na8923_2;
wire na8923_2_i;
wire na8924_1;
wire na8924_1_i;
wire na8924_9;
wire na8925_2;
wire na8925_2_i;
wire na8926_1;
wire na8926_1_i;
wire na8926_9;
wire na8927_2;
wire na8927_2_i;
wire na8928_1;
wire na8928_1_i;
wire na8928_9;
wire na8929_2;
wire na8929_2_i;
wire na8930_1;
wire na8930_1_i;
wire na8930_9;
wire na8931_2;
wire na8931_2_i;
wire na8932_1;
wire na8932_1_i;
wire na8932_9;
wire na8933_2;
wire na8933_2_i;
wire na8934_1;
wire na8934_1_i;
wire na8934_9;
wire na8935_2;
wire na8935_2_i;
wire na8936_1;
wire na8936_1_i;
wire na8936_9;
wire na8937_2;
wire na8937_2_i;
wire na8938_1;
wire na8938_1_i;
wire na8938_9;
wire na8939_2;
wire na8939_2_i;
wire na8940_1;
wire na8940_1_i;
wire na8940_9;
wire na8941_2;
wire na8941_2_i;
wire na8942_1;
wire na8942_1_i;
wire na8942_9;
wire na8943_2;
wire na8943_2_i;
wire na8944_1;
wire na8944_1_i;
wire na8944_9;
wire na8945_2;
wire na8945_2_i;
wire na8946_1;
wire na8946_1_i;
wire na8946_9;
wire na8947_2;
wire na8947_2_i;
wire na8948_1;
wire na8948_1_i;
wire na8948_9;
wire na8949_2;
wire na8950_1;
wire na8950_9;
wire na8951_2;
wire na8952_1;
wire na8952_9;
wire na8953_2;
wire na8954_1;
wire na8954_9;
wire na8955_2;
wire na8956_1;
wire na8956_9;
wire na8957_2;
wire na8958_1;
wire na8958_9;
wire na8959_2;
wire na8960_1;
wire na8960_9;
wire na8961_2;
wire na8962_1;
wire na8962_9;
wire na8963_2;
wire na8964_1;
wire na8964_9;
wire na8965_2;
wire na8966_1;
wire na8966_9;
wire na8967_2;
wire na8968_1;
wire na8968_9;
wire na8969_2;
wire na8970_1;
wire na8970_9;
wire na8971_2;
wire na8972_1;
wire na8972_9;
wire na8973_2;
wire na8974_1;
wire na8974_9;
wire na8975_2;
wire na8976_1;
wire na8976_9;
wire na8977_2;
wire na8978_1;
wire na8978_9;
wire na8979_2;
wire na8980_1;
wire na8980_9;
wire na8981_2;
wire na8982_1;
wire na8982_9;
wire na8983_2;
wire na8984_1;
wire na8984_9;
wire na8985_2;
wire na8986_1;
wire na8986_9;
wire na8987_2;
wire na8988_1;
wire na8988_9;
wire na8989_1;
wire na8989_9;
wire na8990_1;
wire na8990_9;
wire na8991_2;
wire na8992_2;
wire na8993_2;
wire na8994_1;
wire na8994_9;
wire na8995_2;
wire na8996_1;
wire na8996_9;
wire na8997_2;
wire na8998_1;
wire na8998_9;
wire na8999_2;
wire na9000_1;
wire na9000_9;
wire na9001_2;
wire na9002_1;
wire na9002_9;
wire na9003_2;
wire na9004_1;
wire na9004_9;
wire na9005_2;
wire na9006_1;
wire na9006_9;
wire na9007_2;
wire na9008_1;
wire na9008_9;
wire na9009_2;
wire na9010_1;
wire na9010_9;
wire na9011_2;
wire na9012_1;
wire na9012_9;
wire na9013_2;
wire na9014_1;
wire na9014_9;
wire na9015_2;
wire na9016_1;
wire na9016_9;
wire na9017_2;
wire na9018_1;
wire na9018_9;
wire na9019_2;
wire na9020_1;
wire na9020_9;
wire na9021_2;
wire na9022_1;
wire na9022_9;
wire na9023_2;
wire na9024_1;
wire na9024_9;
wire na9025_2;
wire na9026_1;
wire na9026_9;
wire na9027_2;
wire na9028_1;
wire na9028_9;
wire na9029_2;
wire na9030_1;
wire na9030_9;
wire na9031_2;
wire na9032_1;
wire na9032_9;
wire na9033_2;
wire na9034_1;
wire na9034_9;
wire na9035_2;
wire na9036_1;
wire na9036_9;
wire na9037_2;
wire na9038_1;
wire na9038_9;
wire na9039_2;
wire na9040_1;
wire na9040_9;
wire na9041_2;
wire na9042_1;
wire na9042_9;
wire na9043_2;
wire na9044_1;
wire na9044_9;
wire na9045_2;
wire na9046_1;
wire na9046_9;
wire na9047_2;
wire na9048_1;
wire na9048_9;
wire na9049_2;
wire na9050_1;
wire na9050_9;
wire na9051_2;
wire na9052_1;
wire na9052_9;
wire na9053_2;
wire na9054_1;
wire na9054_9;
wire na9055_2;
wire na9056_1;
wire na9056_9;
wire na9057_2;
wire na9058_1;
wire na9058_9;
wire na9059_2;
wire na9060_1;
wire na9060_9;
wire na9061_2;
wire na9062_1;
wire na9062_9;
wire na9063_2;
wire na9064_1;
wire na9064_9;
wire na9065_2;
wire na9066_1;
wire na9066_9;
wire na9067_2;
wire na9068_1;
wire na9068_9;
wire na9069_2;
wire na9070_1;
wire na9070_9;
wire na9071_2;
wire na9072_1;
wire na9072_9;
wire na9073_2;
wire na9074_1;
wire na9074_9;
wire na9075_2;
wire na9076_1;
wire na9076_9;
wire na9077_2;
wire na9078_1;
wire na9078_9;
wire na9079_2;
wire na9080_1;
wire na9080_9;
wire na9081_2;
wire na9082_1;
wire na9082_9;
wire na9083_2;
wire na9084_1;
wire na9084_9;
wire na9085_2;
wire na9086_1;
wire na9086_9;
wire na9087_2;
wire na9088_1;
wire na9088_9;
wire na9089_2;
wire na9090_1;
wire na9090_9;
wire na9091_2;
wire na9092_1;
wire na9092_9;
wire na9093_2;
wire na9094_1;
wire na9094_9;
wire na9095_2;
wire na9096_1;
wire na9096_9;
wire na9097_2;
wire na9098_1;
wire na9098_9;
wire na9099_2;
wire na9100_1;
wire na9100_9;
wire na9101_2;
wire na9102_1;
wire na9102_9;
wire na9103_2;
wire na9104_1;
wire na9104_9;
wire na9105_2;
wire na9106_1;
wire na9106_9;
wire na9107_2;
wire na9108_1;
wire na9108_9;
wire na9109_2;
wire na9110_1;
wire na9110_9;
wire na9111_2;
wire na9112_1;
wire na9112_9;
wire na9113_2;
wire na9114_1;
wire na9114_9;
wire na9115_2;
wire na9116_1;
wire na9116_9;
wire na9117_2;
wire na9118_1;
wire na9119_2;
wire na9120_1;
wire na9121_2;
wire na9122_1;
wire na9123_2;
wire na9124_1;
wire na9125_2;
wire na9126_1;
wire na9127_2;
wire na9128_1;
wire na9129_2;
wire na9130_1;
wire na9131_2;
wire na9132_1;
wire na9133_2;
wire na9134_2;
wire na9135_2;
wire na9136_2;
wire na9137_2;
wire na9138_2;
wire na9139_2;
wire na9140_2;
wire na9141_2;
wire na9142_2;
wire na9143_2;
wire na9144_2;
wire na9145_2;
wire na9146_2;
wire na9147_2;
wire na9148_2;
wire na9149_2;
wire na9150_2;
wire na9151_2;
wire na9152_2;
wire na9153_2;
wire na9154_2;
wire na9155_2;
wire na9156_2;
wire na9157_2;
wire na9158_2;
wire na9159_2;
wire na9160_2;
wire na9161_2;
wire na9162_2;
wire na9163_2;
wire na9164_2;
wire na9165_2;
wire na9166_2;
wire na9167_2;
wire na9168_2;
wire na9169_2;
wire na9170_2;
wire na9171_2;
wire na9172_2;
wire na9173_2;
wire na9174_2;
wire na9175_2;
wire na9176_2;
wire na9177_2;
wire na9178_2;
wire na9179_2;
wire na9180_2;
wire na9181_2;
wire na9182_2;
wire na9183_2;
wire na9184_2;
wire na9185_2;
wire na9186_2;
wire na9187_2;
wire na9188_2;
wire na9189_2;
wire na9190_2;
wire na9191_2;
wire na9192_2;
wire na9193_2;
wire na9194_2;
wire na9195_2;
wire na9196_2;
wire na9197_2;
wire na9198_2;
wire na9199_2;
wire na9200_2;
wire na9201_2;
wire na9202_2;
wire na9203_2;
wire na9204_2;
wire na9205_2;
wire na9206_2;
wire na9207_2;
wire na9208_2;
wire na9209_2;
wire na9210_2;
wire na9211_2;
wire na9212_2;
wire na9213_2;
wire na9214_2;
wire na9215_2;
wire na9216_2;
wire na9217_2;
wire na9218_2;
wire na9219_2;
wire na9220_2;
wire na9221_2;
wire na9222_2;
wire na9223_2;
wire na9224_2;
wire na9225_2;
wire na9226_2;
wire na9227_2;
wire na9228_2;
wire na9229_2;
wire na9230_2;
wire na9231_2;
wire na9232_2;
wire na9233_2;
wire na9234_2;
wire na9235_2;
wire na9236_2;
wire na9237_2;
wire na9238_2;
wire na9239_2;
wire na9240_2;
wire na9241_2;
wire na9242_2;
wire na9243_2;
wire na9244_2;
wire na9245_2;
wire na9246_2;
wire na9247_2;
wire na9248_2;
wire na9249_2;
wire na9250_2;
wire na9251_2;
wire na9252_2;
wire na9253_2;
wire na9254_2;
wire na9255_2;
wire na9256_2;
wire na9257_2;
wire na9258_2;
wire na9259_2;
wire na9260_2;
wire na9261_2;
wire na9262_2;
wire na9263_2;
wire na9264_2;
wire na9265_2;
wire na9266_2;
wire na9267_2;
wire na9268_2;
wire na9269_2;
wire na9270_2;
wire na9271_2;
wire na9272_2;
wire na9273_2;
wire na9274_2;
wire na9275_2;
wire na9276_2;
wire na9277_2;
wire na9278_2;
wire na9279_2;
wire na9280_2;
wire na9281_2;
wire na9282_2;
wire na9283_2;
wire na9284_2;
wire na9285_2;
wire na9286_2;
wire na9287_2;
wire na9288_2;
wire na9289_2;
wire na9290_2;
wire na9291_2;
wire na9292_2;
wire na9293_2;
wire na9294_2;
wire na9295_2;
wire na9296_2;
wire na9297_2;
wire na9298_2;
wire na9299_2;
wire na9300_2;
wire na9301_2;
wire na9302_2;
wire na9303_2;
wire na9304_2;
wire na9305_2;
wire na9306_2;
wire na9307_2;
wire na9308_2;
wire na9309_2;
wire na9310_2;
wire na9311_2;
wire na9312_2;
wire na9313_2;
wire na9314_2;
wire na9315_2;
wire na9316_2;
wire na9317_2;
wire na9318_2;
wire na9319_2;
wire na9320_2;
wire na9321_2;
wire na9322_2;
wire na9323_2;
wire na9324_2;
wire na9325_2;
wire na9326_2;
wire na9327_2;
wire na9328_2;
wire na9329_2;
wire na9330_2;
wire na9331_2;
wire na9332_2;
wire na9333_2;
wire na9334_2;
wire na9335_2;
wire na9336_2;
wire na9337_2;
wire na9338_2;
wire na9339_2;
wire na9340_2;
wire na9341_2;
wire na9342_2;
wire na9343_2;
wire na9344_2;
wire na9345_2;
wire na9346_2;
wire na9347_2;
wire na9348_2;
wire na9349_2;
wire na9350_2;
wire na9351_2;
wire na9352_2;
wire na9353_2;
wire na9354_2;
wire na9355_2;
wire na9356_2;
wire na9357_2;
wire na9358_2;
wire na9359_2;
wire na9360_2;
wire na9361_2;
wire na9362_2;
wire na9363_2;
wire na9364_2;
wire na9365_2;
wire na9366_2;
wire na9367_2;
wire na9368_2;
wire na9369_2;
wire na9370_2;
wire na9371_2;
wire na9372_2;
wire na9373_2;
wire na9374_2;
wire na9375_2;
wire na9376_2;
wire na9377_2;
wire na9378_2;
wire na9379_2;
wire na9380_2;
wire na9381_2;
wire na9382_2;
wire na9383_2;
wire na9384_2;
wire na9385_2;
wire na9386_2;
wire na9387_2;
wire na9388_2;
wire na9389_2;
wire na9390_2;
wire na9391_2;
wire na9392_2;
wire na9393_2;
wire na9394_2;
wire na9395_2;
wire na9396_2;
wire na9397_2;
wire na9398_2;
wire na9399_2;
wire na9400_2;
wire na9401_2;
wire na9402_2;
wire na9403_2;
wire na9404_2;
wire na9405_2;
wire na9406_2;
wire na9407_2;
wire na9408_2;
wire na9409_2;
wire na9410_2;
wire na9411_2;
wire na9412_2;
wire na9413_2;
wire na9414_2;
wire na9415_2;
wire na9416_2;
wire na9417_2;
wire na9418_2;
wire na9419_2;
wire na9420_2;
wire na9421_2;
wire na9422_2;
wire na9423_2;
wire na9424_2;
wire na9425_2;
wire na9426_2;
wire na9427_2;
wire na9428_2;
wire na9429_2;
wire na9430_2;
wire na9431_2;
wire na9432_2;
wire na9433_2;
wire na9434_2;
wire na9435_2;
wire na9436_2;
wire na9437_2;
wire na9438_2;
wire na9439_2;
wire na9440_2;
wire na9441_2;
wire na9442_2;
wire na9443_2;
wire na9444_2;
wire na9445_2;
wire na9446_2;
wire na9447_2;
wire na9448_2;
wire na9449_2;
wire na9450_2;
wire na9451_2;
wire na9452_2;
wire na9453_2;
wire na9454_2;
wire na9455_2;
wire na9456_2;
wire na9457_2;
wire na9458_2;
wire na9459_2;
wire na9460_2;
wire na9461_2;
wire na9462_2;
wire na9463_2;
wire na9464_2;
wire na9465_2;
wire na9466_2;
wire na9467_2;
wire na9468_2;
wire na9469_2;
wire na9470_2;
wire na9471_2;
wire na9472_2;
wire na9473_2;
wire na9474_2;
wire na9475_2;
wire na9476_2;
wire na9477_2;
wire na9478_2;
wire na9479_2;
wire na9480_2;
wire na9481_2;
wire na9482_2;
wire na9483_2;
wire na9484_2;
wire na9485_2;
wire na9486_2;
wire na9487_2;
wire na9488_2;
wire na9489_2;
wire na9490_2;
wire na9491_2;
wire na9492_2;
wire na9493_2;
wire na9494_2;
wire na9495_2;
wire na9496_2;
wire na9497_2;
wire na9498_2;
wire na9499_2;
wire na9500_2;
wire na9501_2;
wire na9502_2;
wire na9503_2;
wire na9504_2;
wire na9505_2;
wire na9506_2;
wire na9507_2;
wire na9508_2;
wire na9509_2;
wire na9510_2;
wire na9511_2;
wire na9512_2;
wire na9513_2;
wire na9514_2;
wire na9515_2;
wire na9516_2;
wire na9517_2;
wire na9518_2;
wire na9519_2;
wire na9520_2;
wire na9521_2;
wire na9522_2;
wire na9523_2;
wire na9524_2;
wire na9525_2;
wire na9526_2;
wire na9527_2;
wire na9528_2;
wire na9529_2;
wire na9530_2;
wire na9531_2;
wire na9532_2;
wire na9533_2;
wire na9534_2;
wire na9535_2;
wire na9536_2;
wire na9537_2;
wire na9538_2;
wire na9539_2;
wire na9540_2;
wire na9541_2;
wire na9542_2;
wire na9543_2;
wire na9544_2;
wire na9545_2;
wire na9546_2;
wire na9547_2;
wire na9548_2;
wire na9549_2;
wire na9550_2;
wire na9551_2;
wire na9552_2;
wire na9553_2;
wire na9554_2;
wire na9555_2;
wire na9556_2;
wire na9557_2;
wire na9558_2;
wire na9559_2;
wire na9560_2;
wire na9561_2;
wire na9562_2;
wire na9563_2;
wire na9564_2;
wire na9565_2;
wire na9566_2;
wire na9567_2;
wire na9568_2;
wire na9569_2;
wire na9570_2;
wire na9571_2;
wire na9572_2;
wire na9573_2;
wire na9574_2;
wire na9575_2;
wire na9576_2;
wire na9577_2;
wire na9578_2;
wire na9579_2;
wire na9580_2;
wire na9581_2;
wire na9582_2;
wire na9583_2;
wire na9584_2;
wire na9585_2;
wire na9586_2;
wire na9587_2;
wire na9588_2;
wire na9589_2;
wire na9590_2;
wire na9591_2;
wire na9592_2;
wire na9593_2;
wire na9594_2;
wire na9595_2;
wire na9596_2;
wire na9597_2;
wire na9598_2;
wire na9599_2;
wire na9600_2;
wire na9601_2;
wire na9602_2;
wire na9603_2;
wire na9604_2;
wire na9605_2;
wire na9606_2;
wire na9607_2;
wire na9608_2;
wire na9609_2;
wire na9610_2;
wire na9611_2;
wire na9612_2;
wire na9613_2;
wire na9614_2;
wire na9615_2;
wire na9616_2;
wire na9617_2;
wire na9618_2;
wire na9619_2;
wire na9620_2;
wire na9621_2;
wire na9622_2;
wire na9623_2;
wire na9624_2;
wire na9625_2;
wire na9626_2;
wire na9627_2;
wire na9628_2;
wire na9629_2;
wire na9630_2;
wire na9631_2;
wire na9632_2;
wire na9633_2;
wire na9634_2;
wire na9635_2;
wire na9636_2;
wire na9637_2;
wire na9638_2;
wire na9639_2;
wire na9640_2;
wire na9641_2;
wire na9642_2;
wire na9643_2;
wire na9644_2;
wire na9645_2;
wire na9646_2;
wire na9647_2;
wire na9648_2;
wire na9649_2;
wire na9650_2;
wire na9651_2;
wire na9652_2;
wire na9653_2;
wire na9654_2;
wire na9655_2;
wire na9656_2;
wire na9657_2;
wire na9658_2;
wire na9659_2;
wire na9660_2;
wire na9661_2;
wire na9662_2;
wire na9663_2;
wire na9664_2;
wire na9665_2;
wire na9666_2;
wire na9667_2;
wire na9668_2;
wire na9669_2;
wire na9670_2;
wire na9671_2;
wire na9672_2;
wire na9673_2;
wire na9674_2;
wire na9675_2;
wire na9676_2;
wire na9677_2;
wire na9678_2;
wire na9679_2;
wire na9680_2;
wire na9681_2;
wire na9682_2;
wire na9683_2;
wire na9684_2;
wire na9685_2;
wire na9686_2;
wire na9687_2;
wire na9688_2;
wire na9689_2;
wire na9690_2;
wire na9691_2;
wire na9692_2;
wire na9693_2;
wire na9694_2;
wire na9695_2;
wire na9696_2;
wire na9697_2;
wire na9698_2;
wire na9699_2;
wire na9700_2;
wire na9701_2;
wire na9702_2;
wire na9703_2;
wire na9704_2;
wire na9705_2;
wire na9706_2;
wire na9707_2;
wire na9708_2;
wire na9709_2;
wire na9710_2;
wire na9711_2;
wire na9712_2;
wire na9713_2;
wire na9714_2;
wire na9715_2;
wire na9716_2;
wire na9717_2;
wire na9718_2;
wire na9719_2;
wire na9720_2;
wire na9721_2;
wire na9722_2;
wire na9723_2;
wire na9724_2;
wire na9725_2;
wire na9726_2;
wire na9727_2;
wire na9728_2;
wire na9729_2;
wire na9730_2;
wire na9731_2;
wire na9732_2;
wire na9733_2;
wire na9734_2;
wire na9735_2;
wire na9736_2;
wire na9737_2;
wire na9738_2;
wire na9739_2;
wire na9740_2;
wire na9741_2;
wire na9742_2;
wire na9743_2;
wire na9744_2;
wire na9745_2;
wire na9746_2;
wire na9747_2;
wire na9748_2;
wire na9749_2;
wire na9750_2;
wire na9751_2;
wire na9752_2;
wire na9753_2;
wire na9754_2;
wire na9755_2;
wire na9756_2;
wire na9757_2;
wire na9758_2;
wire na9759_2;
wire na9760_2;
wire na9761_2;
wire na9762_2;
wire na9763_2;
wire na9764_2;
wire na9765_2;
wire na9766_2;
wire na9767_2;
wire na9768_2;
wire na9769_2;
wire na9770_2;
wire na9771_2;
wire na9772_2;
wire na9773_2;
wire na9774_2;
wire na9775_2;
wire na9776_2;
wire na9777_2;
wire na9778_2;
wire na9779_2;
wire na9780_2;
wire na9781_2;
wire na9782_2;
wire na9783_2;
wire na9784_2;
wire na9785_2;
wire na9786_2;
wire na9787_2;
wire na9788_2;
wire na9789_2;
wire na9790_2;
wire na9791_2;
wire na9792_2;
wire na9793_2;
wire na9794_2;
wire na9795_2;
wire na9796_2;
wire na9797_2;
wire na9798_2;
wire na9799_2;
wire na9800_2;
wire na9801_2;
wire na9802_2;
wire na9803_2;
wire na9804_2;
wire na9805_2;
wire na9806_2;
wire na9807_2;
wire na9808_2;
wire na9809_2;
wire na9810_2;
wire na9811_2;
wire na9812_2;
wire na9813_2;
wire na9814_2;
wire na9815_2;
wire na9816_2;
wire na9817_2;
wire na9818_2;
wire na9819_2;
wire na9820_2;
wire na9821_2;
wire na9822_2;
wire na9823_2;
wire na9824_2;
wire na9825_2;
wire na9826_2;
wire na9827_2;
wire na9828_2;
wire na9829_2;
wire na9830_2;
wire na9831_2;
wire na9832_2;
wire na9833_2;
wire na9834_2;
wire na9835_2;
wire na9836_2;
wire na9837_2;
wire na9838_2;
wire na9839_2;
wire na9840_2;
wire na9841_2;
wire na9842_2;
wire na9843_2;
wire na9844_2;
wire na9845_2;
wire na9846_2;
wire na9847_2;
wire na9848_2;
wire na9849_2;
wire na9850_2;
wire na9851_2;
wire na9852_2;
wire na9853_2;
wire na9854_2;
wire na9855_2;
wire na9856_2;
wire na9857_2;
wire na9858_2;
wire na9859_2;
wire na9860_2;
wire na9861_2;
wire na9862_2;
wire na9863_2;
wire na9864_2;
wire na9865_2;
wire na9866_2;
wire na9867_2;
wire na9868_2;
wire na9869_2;
wire na9870_2;
wire na9871_2;
wire na9872_2;
wire na9873_2;
wire na9874_2;
wire na9875_2;
wire na9876_2;
wire na9877_2;
wire na9878_2;
wire na9879_2;
wire na9880_2;
wire na9881_2;
wire na9882_2;
wire na9883_2;
wire na9884_2;
wire na9885_2;
wire na9886_2;
wire na9887_2;
wire na9888_2;
wire na9889_2;
wire na9890_2;
wire na9891_2;
wire na9892_2;
wire na9893_2;
wire na9894_2;
wire na9895_2;
wire na9896_2;
wire na9897_2;
wire na9898_2;
wire na9899_2;
wire na9900_2;
wire na9901_2;
wire na9902_2;
wire na9903_2;
wire na9904_2;
wire na9905_2;
wire na9906_2;
wire na9907_2;
wire na9908_2;
wire na9909_2;
wire na9910_2;
wire na9911_2;
wire na9912_2;
wire na9913_2;
wire na9914_2;
wire na9915_2;
wire na9916_2;
wire na9917_2;
wire na9918_2;
wire na9919_2;
wire na9920_2;
wire na9921_2;
wire na9922_2;
wire na9923_2;
wire na9924_2;
wire na9925_2;
wire na9926_2;
wire na9927_2;
wire na9928_2;
wire na9929_2;
wire na9930_2;
wire na9931_2;
wire na9932_2;
wire na9933_2;
wire na9934_2;
wire na9935_2;
wire na9936_2;
wire na9937_2;
wire na9938_2;
wire na9939_2;
wire na9940_2;
wire na9941_2;
wire na9942_2;
wire na9943_2;
wire na9944_2;
wire na9945_2;
wire na9946_2;
wire na9947_2;
wire na9948_2;
wire na9949_2;
wire na9950_2;
wire na9951_2;
wire na9952_2;
wire na9953_2;
wire na9954_2;
wire na9955_2;
wire na9956_2;
wire na9957_2;
wire na9958_2;
wire na9959_2;
wire na9960_2;
wire na9961_2;
wire na9962_2;
wire na9963_2;
wire na9964_2;
wire na9965_2;
wire na9966_2;
wire na9967_2;
wire na9968_2;
wire na9969_2;
wire na9970_2;
wire na9971_2;
wire na9972_2;
wire na9973_2;
wire na9974_2;
wire na9975_2;
wire na9976_2;
wire na9977_2;
wire na9978_2;
wire na9979_2;
wire na9980_2;
wire na9981_2;
wire na9982_2;
wire na9983_2;
wire na9984_2;
wire na9985_2;
wire na9986_2;
wire na9987_2;
wire na9988_2;
wire na9989_2;
wire na9990_2;
wire na9991_2;
wire na9992_2;
wire na9993_2;
wire na9994_2;
wire na9995_2;
wire na9996_2;
wire na9997_2;
wire na9998_2;
wire na9999_2;
wire cdone_ice40;
wire na10000_2;
wire na10001_2;
wire na10002_2;
wire na10003_2;
wire na10004_2;
wire na10005_2;
wire na10006_2;
wire na10007_2;
wire na10008_2;
wire na10009_2;
wire na10010_2;
wire na10011_2;
wire na10012_2;
wire na10013_2;
wire na10014_2;
wire na10015_2;
wire na10016_2;
wire na10017_2;
wire na10018_2;
wire na10019_2;
wire na10020_2;
wire na10021_2;
wire na10022_2;
wire na10023_2;
wire na10024_2;
wire na10025_2;
wire na10026_2;
wire na10027_2;
wire na10028_2;
wire na10029_2;
wire na10030_2;
wire na10031_2;
wire na10032_2;
wire na10033_2;
wire na10034_2;
wire na10035_2;
wire na10036_2;
wire na10037_2;
wire na10038_2;
wire na10039_2;
wire na10040_2;
wire na10041_2;
wire na10042_2;
wire na10043_2;
wire na10044_2;
wire na10045_2;
wire na10046_2;
wire na10047_2;
wire na10048_2;
wire na10049_2;
wire na10050_2;
wire na10051_2;
wire na10052_2;
wire na10053_2;
wire na10054_2;
wire na10055_2;
wire na10056_2;
wire na10057_2;
wire na10058_2;
wire na10059_2;
wire na10060_2;
wire na10061_2;
wire na10062_2;
wire na10063_2;
wire na10064_2;
wire na10065_2;
wire na10066_2;
wire na10067_2;
wire na10068_2;
wire na10069_2;
wire na10070_2;
wire na10071_2;
wire na10072_2;
wire na10073_2;
wire na10074_2;
wire na10075_2;
wire na10076_2;
wire na10077_2;
wire na10078_2;
wire na10079_2;
wire na10080_2;
wire na10081_2;
wire na10082_2;
wire na10083_2;
wire na10084_2;
wire na10085_2;
wire na10086_2;
wire na10087_2;
wire na10088_2;
wire na10089_2;
wire na10090_2;
wire na10091_2;
wire na10092_2;
wire na10093_2;
wire na10094_2;
wire na10095_2;
wire na10096_2;
wire na10097_2;
wire na10098_2;
wire na10099_2;
wire na10100_2;
wire na10101_2;
wire na10102_2;
wire na10103_2;
wire na10104_2;
wire na10105_2;
wire na10106_2;
wire na10107_2;
wire na10108_2;
wire na10109_2;
wire na10110_2;
wire na10111_2;
wire na10112_2;
wire na10113_2;
wire na10114_2;
wire na10115_2;
wire na10116_2;
wire na10117_2;
wire na10118_2;
wire na10119_2;
wire na10120_2;
wire na10121_2;
wire na10122_2;
wire na10123_2;
wire na10124_2;
wire na10125_2;
wire na10126_2;
wire na10127_2;
wire na10128_2;
wire na10129_2;
wire na10130_2;
wire na10131_2;
wire na10132_2;
wire na10133_2;
wire na10134_2;
wire na10135_2;
wire na10136_2;
wire na10137_2;
wire na10138_2;
wire na10139_2;
wire na10140_2;
wire na10141_2;
wire na10142_2;
wire na10143_2;
wire na10144_2;
wire na10145_2;
wire na10146_2;
wire na10147_2;
wire na10148_2;
wire na10149_2;
wire na10150_2;
wire na10151_2;
wire na10152_2;
wire na10153_2;
wire na10154_2;
wire na10155_2;
wire na10156_2;
wire na10157_2;
wire na10158_2;
wire na10159_2;
wire na10160_2;
wire na10161_2;
wire na10162_2;
wire na10163_2;
wire na10164_2;
wire na6629_21;
wire na6629_22;
wire na6629_23;
wire na6629_24;
wire na6629_25;
wire na6629_26;
wire na6629_27;
wire na6629_28;
wire na6629_29;
wire na6629_30;
wire na6629_31;
wire na6629_32;
wire na6629_33;
wire na6629_34;
wire na6629_35;
wire na6629_36;
wire na6629_37;
wire na6629_38;
wire na6629_39;
wire na6629_40;
wire na6630_10;
wire na6630_11;
wire na6630_12;
wire na6630_13;
wire na6630_14;
wire na6630_15;
wire na6630_16;
wire na6630_17;
wire na6630_18;
wire na6630_19;
wire na6630_20;
wire na6630_89;
wire na6630_90;
wire na6630_91;
wire na6630_92;
wire na6630_93;
wire na6630_94;
wire na6630_95;
wire na6630_96;
wire na6630_97;
wire na6630_98;
wire na6630_99;
wire na6631_36;
wire na6631_37;
wire na6631_38;
wire na6631_39;
wire na6631_40;
wire na6632_36;
wire na6632_37;
wire na6632_38;
wire na6632_39;
wire na6632_40;
wire na6633_36;
wire na6633_37;
wire na6633_38;
wire na6633_39;
wire na6633_40;
wire na6634_36;
wire na6634_37;
wire na6634_38;
wire na6634_39;
wire na6634_40;
wire na6635_37;
wire na6635_38;
wire na6635_39;
wire na6635_40;
wire na6636_36;
wire na6636_37;
wire na6636_38;
wire na6636_39;
wire na6636_40;
wire na6637_36;
wire na6637_37;
wire na6637_38;
wire na6637_39;
wire na6637_40;
wire na6638_36;
wire na6638_37;
wire na6638_38;
wire na6638_39;
wire na6638_40;
wire na6639_36;
wire na6639_37;
wire na6639_38;
wire na6639_39;
wire na6639_40;
wire na6640_36;
wire na6640_37;
wire na6640_38;
wire na6640_39;
wire na6640_40;
wire na6641_36;
wire na6641_37;
wire na6641_38;
wire na6641_39;
wire na6641_40;
wire na6642_36;
wire na6642_37;
wire na6642_38;
wire na6642_39;
wire na6642_40;
wire na6643_36;
wire na6643_37;
wire na6643_38;
wire na6643_39;
wire na6643_40;
wire na6644_21;
wire na6644_22;
wire na6644_23;
wire na6644_24;
wire na6644_25;
wire na6644_26;
wire na6644_27;
wire na6644_28;
wire na6644_29;
wire na6644_30;
wire na6644_31;
wire na6644_32;
wire na6644_33;
wire na6644_34;
wire na6644_35;
wire na6644_36;
wire na6644_37;
wire na6644_38;
wire na6644_39;
wire na6644_40;
wire na6645_10;
wire na6645_11;
wire na6645_12;
wire na6645_13;
wire na6645_14;
wire na6645_15;
wire na6645_16;
wire na6645_17;
wire na6645_18;
wire na6645_19;
wire na6645_20;
wire na6645_21;
wire na6645_22;
wire na6645_23;
wire na6645_24;
wire na6645_25;
wire na6645_26;
wire na6645_27;
wire na6645_28;
wire na6645_29;
wire na6645_30;
wire na6645_31;
wire na6645_32;
wire na6645_33;
wire na6645_34;
wire na6645_35;
wire na6645_36;
wire na6645_37;
wire na6645_38;
wire na6645_39;
wire na6645_40;
wire na6646_10;
wire na6647_21;
wire na6647_22;
wire na6647_23;
wire na6647_24;
wire na6647_25;
wire na6647_26;
wire na6647_27;
wire na6647_28;
wire na6647_29;
wire na6647_30;
wire na6647_31;
wire na6647_32;
wire na6647_33;
wire na6647_34;
wire na6647_35;
wire na6647_36;
wire na6647_37;
wire na6647_38;
wire na6647_39;
wire na6647_40;
wire na6648_10;
wire na6648_11;
wire na6648_12;
wire na6648_13;
wire na6648_14;
wire na6648_15;
wire na6648_16;
wire na6648_17;
wire na6648_18;
wire na6648_19;
wire na6648_20;
wire na6648_21;
wire na6648_22;
wire na6648_23;
wire na6648_24;
wire na6648_25;
wire na6648_26;
wire na6648_27;
wire na6648_28;
wire na6648_29;
wire na6648_30;
wire na6648_31;
wire na6648_32;
wire na6648_33;
wire na6648_34;
wire na6648_35;
wire na6648_36;
wire na6648_37;
wire na6648_38;
wire na6648_39;
wire na6648_40;
wire na6649_10;
wire na6650_10;
wire na6650_11;
wire na6650_12;
wire na6650_13;
wire na6650_14;
wire na6650_15;
wire na6650_16;
wire na6650_17;
wire na6650_18;
wire na6650_19;
wire na6650_20;
wire na6650_33;
wire na6650_34;
wire na6650_35;
wire na6650_36;
wire na6650_37;
wire na6650_38;
wire na6650_39;
wire na6650_40;
wire na6651_10;
wire na6651_11;
wire na6651_12;
wire na6651_13;
wire na6651_14;
wire na6651_15;
wire na6651_16;
wire na6651_17;
wire na6651_18;
wire na6651_19;
wire na6651_20;
wire na6651_21;
wire na6651_22;
wire na6651_23;
wire na6651_24;
wire na6651_25;
wire na6651_26;
wire na6651_27;
wire na6651_28;
wire na6651_29;
wire na6651_30;
wire na6651_31;
wire na6651_32;
wire na6651_33;
wire na6651_34;
wire na6651_35;
wire na6651_36;
wire na6651_37;
wire na6651_38;
wire na6651_39;
wire na6651_40;
wire na6653_10;
wire na6653_11;
wire na6653_12;
wire na6653_13;
wire na6653_14;
wire na6653_15;
wire na6653_16;
wire na6653_17;
wire na6653_18;
wire na6653_19;
wire na6653_20;
wire na6653_21;
wire na6653_22;
wire na6653_23;
wire na6653_24;
wire na6653_25;
wire na6653_26;
wire na6653_27;
wire na6653_28;
wire na6653_29;
wire na6653_30;
wire na6653_31;
wire na6653_32;
wire na6653_33;
wire na6653_34;
wire na6653_35;
wire na6653_36;
wire na6653_37;
wire na6653_38;
wire na6653_39;
wire na6653_40;
wire na6654_10;
wire na6655_21;
wire na6655_22;
wire na6655_23;
wire na6655_24;
wire na6655_25;
wire na6655_26;
wire na6655_27;
wire na6655_28;
wire na6655_29;
wire na6655_30;
wire na6655_31;
wire na6655_32;
wire na6655_33;
wire na6655_34;
wire na6655_35;
wire na6655_36;
wire na6655_37;
wire na6655_38;
wire na6655_39;
wire na6655_40;
wire na6657_10;
wire na6657_11;
wire na6657_12;
wire na6657_13;
wire na6657_14;
wire na6657_15;
wire na6657_16;
wire na6657_17;
wire na6657_18;
wire na6657_19;
wire na6657_20;
wire na6657_21;
wire na6657_22;
wire na6657_23;
wire na6657_24;
wire na6657_25;
wire na6657_26;
wire na6657_27;
wire na6657_28;
wire na6657_29;
wire na6657_30;
wire na6657_31;
wire na6657_32;
wire na6657_33;
wire na6657_34;
wire na6657_35;
wire na6657_36;
wire na6657_37;
wire na6657_38;
wire na6657_39;
wire na6657_40;
wire na6658_10;
wire na6659_93;
wire na6659_94;
wire na6659_95;
wire na6659_96;
wire na6659_97;
wire na6659_98;
wire na6659_99;
wire na6667_10;
wire na6670_10;
wire na6679_10;
wire na6682_10;
wire na6685_10;
wire na6687_10;
wire na6689_10;
wire na6691_10;
wire na6694_10;
wire na6698_10;
wire na6704_10;
wire na6708_10;
wire na6714_10;
wire na6716_10;
wire na6718_10;
wire na6721_10;
wire na6725_10;
wire na6728_10;
wire na6730_10;
wire na6732_10;
wire na6735_10;
wire na6738_10;
wire na6740_10;
wire na6744_10;
wire na6747_10;
wire na6751_10;
wire na6755_10;
wire na6757_10;
wire na6760_10;
wire na6762_10;
wire na6764_10;
wire na6766_10;
wire na6773_10;
wire na6791_10;
wire na6793_10;
wire na6800_10;
wire na6802_10;
wire na6806_10;
wire na6809_10;
wire na6813_10;
wire na6815_10;
wire na6818_10;
wire na6820_10;
wire na6822_10;
wire na6825_10;
wire na6827_10;
wire na6830_10;
wire na6832_10;
wire na6835_10;
wire na6838_10;
wire na6842_10;
wire na6844_10;
wire na6848_10;
wire na6851_10;
wire na6854_10;
wire na6857_10;
wire na6860_10;
wire na6862_10;
wire na6865_10;
wire na6873_10;
wire na6876_10;
wire na6878_10;
wire na6882_10;
wire na6884_10;
wire na6890_10;
wire na6894_10;
wire na6897_10;
wire na6899_10;
wire na6902_10;
wire na6905_10;
wire na6908_10;
wire na6911_10;
wire na6914_10;
wire na6916_10;
wire na6919_10;
wire na6922_10;
wire na6924_10;
wire na6927_10;
wire na6930_10;
wire na6932_10;
wire na6939_10;
wire na6949_10;
wire na6952_10;
wire na6955_10;
wire na6957_10;
wire na6960_10;
wire na6963_10;
wire na6965_10;
wire na6968_10;
wire na6971_10;
wire na6973_10;
wire na6976_10;
wire na6986_10;
wire na6989_10;
wire na6993_10;
wire na7000_10;
wire na7005_10;
wire na7013_10;
wire na7030_10;
wire na7037_10;
wire na7048_10;
wire na7053_10;
wire na7058_10;
wire na7070_10;
wire na7074_10;
wire na7077_10;
wire na7080_10;
wire na7083_10;
wire na7085_10;
wire na7088_10;
wire na7091_10;
wire na7093_10;
wire na7099_10;
wire na7103_10;
wire na7116_10;
wire na7119_10;
wire na7123_10;
wire na7126_10;
wire na7128_10;
wire na7137_10;
wire na7139_10;
wire na7149_10;
wire na7151_10;
wire na7155_10;
wire na7159_10;
wire na7169_10;
wire na7172_10;
wire na7174_10;
wire na7177_10;
wire na7180_10;
wire na7193_10;
wire na7195_10;
wire na7197_10;
wire na7200_10;
wire na7205_10;
wire na7214_10;
wire na7225_10;
wire na7227_10;
wire na7230_10;
wire na7236_10;
wire na7238_10;
wire na7241_10;
wire na7243_10;
wire na7246_10;
wire na7248_10;
wire na7251_10;
wire na7253_10;
wire na7267_10;
wire na7269_10;
wire na7272_10;
wire na7274_10;
wire na7280_10;
wire na7284_10;
wire na7287_10;
wire na7289_10;
wire na7303_10;
wire na7306_10;
wire na7308_10;
wire na7331_10;
wire na7333_10;
wire na7337_10;
wire na7340_10;
wire na7342_10;
wire na7350_10;
wire na7352_10;
wire na7356_10;
wire na7358_10;
wire na7365_10;
wire na7368_10;
wire na7379_10;
wire na7382_10;
wire na7384_10;
wire na7387_10;
wire na7390_10;
wire na7392_10;
wire na7395_10;
wire na7398_10;
wire na7400_10;
wire na7403_10;
wire na7406_10;
wire na7416_10;
wire na7419_10;
wire na7422_10;
wire na7424_10;
wire na7427_10;
wire na7430_10;
wire na7432_10;
wire na7435_10;
wire na7438_10;
wire na7440_10;
wire na7443_10;
wire na7454_10;
wire na7456_10;
wire na7459_10;
wire na7462_10;
wire na7464_10;
wire na7467_10;
wire na7470_10;
wire na7472_10;
wire na7475_10;
wire na7478_10;
wire na7480_10;
wire na7499_10;
wire na7502_10;
wire na7504_10;
wire na7507_10;
wire na7510_10;
wire na7512_10;
wire na7515_10;
wire na7518_10;
wire na7520_10;
wire na7523_10;
wire na7526_10;
wire na7536_10;
wire na7538_10;
wire na7540_10;
wire na7543_10;
wire na7546_10;
wire na7548_10;
wire na7551_10;
wire na7554_10;
wire na7556_10;
wire na7562_10;
wire na7564_10;
wire na7567_10;
wire na7570_10;
wire na7572_10;
wire na7575_10;
wire na7578_10;
wire na7580_10;
wire na7583_10;
wire na7586_10;
wire na7588_10;
wire na7591_10;
wire na7602_10;
wire na7604_10;
wire na7607_10;
wire na7618_10;
wire na7620_10;
wire na7625_10;
wire na7631_10;
wire na7635_10;
wire na7638_10;
wire na7640_10;
wire na7646_10;
wire na7647_10;
wire na7648_10;
wire na7651_10;
wire na7654_10;
wire na7656_10;
wire na7659_10;
wire na7710_10;
wire na7712_10;
wire na7715_10;
wire na7717_10;
wire na7719_10;
wire na7721_10;
wire na7724_10;
wire na7726_10;
wire na7734_10;
wire na7742_10;
wire na7750_10;
wire na7766_10;
wire na7777_10;
wire na7789_10;
wire na7795_10;
wire na7801_10;
wire na7807_10;
wire na7813_10;
wire na7819_10;
wire na7827_10;
wire na7835_10;
wire na7843_10;
wire na7851_10;
wire na7859_10;
wire na7867_10;
wire na7875_10;
wire na7883_10;
wire na7892_10;
wire na7896_10;
wire na7900_10;
wire na7904_10;
wire na7907_10;
wire na7909_10;
wire na7913_10;
wire na7915_10;
wire na7917_10;
wire na7920_10;
wire na7923_10;
wire na7927_10;
wire na7931_10;
wire na7933_10;
wire na7937_10;
wire na7941_10;
wire na7945_10;
wire na7947_10;
wire na7951_10;
wire na7958_10;
wire na7962_10;
wire na7965_10;
wire na7969_10;
wire na7972_10;
wire na7974_10;
wire na7977_10;
wire na7980_10;
wire na7982_10;
wire na7986_10;
wire na7988_10;
wire na7990_10;
wire na7992_10;
wire na7995_10;
wire na7998_10;
wire na8001_10;
wire na8004_10;
wire na8007_10;
wire na8013_10;
wire na8016_10;
wire na8019_10;
wire na8022_10;
wire na8025_10;
wire na8028_10;
wire na8031_10;
wire na8034_10;
wire na8037_10;
wire na8040_10;
wire na8042_10;
wire na8044_10;
wire na8046_10;
wire na8048_10;
wire na8050_10;
wire na8052_10;
wire na8054_10;
wire na8056_10;
wire na8059_10;
wire na8062_10;
wire na8066_10;
wire na8071_10;
wire na8083_10;
wire na8084_10;
wire na8086_10;
wire na8090_10;
wire na8102_10;
wire na8108_10;
wire na8112_10;
wire na8115_10;
wire na8120_10;
wire na8124_10;
wire na8127_10;
wire na8129_10;
wire na8133_10;
wire na8136_10;
wire na8139_10;
wire na8141_10;
wire na8144_10;
wire na8146_10;
wire na8150_10;
wire na8155_10;
wire na8160_10;
wire na8162_10;
wire na8164_10;
wire na8168_10;
wire na8170_10;
wire na8172_10;
wire na8179_10;
wire na8181_10;
wire na8189_10;
wire na8193_10;
wire na8195_10;
wire na8198_10;
wire na8200_10;
wire na8202_10;
wire na8204_10;
wire na8206_10;
wire na8208_10;
wire na8210_10;
wire na8212_10;
wire na8214_10;
wire na8216_10;
wire na8218_10;
wire na8220_10;
wire na8222_10;
wire na8224_10;
wire na8226_10;
wire na8228_10;
wire na8230_10;
wire na8232_10;
wire na8234_10;
wire na8236_10;
wire na8238_10;
wire na8240_10;
wire na8242_10;
wire na8244_10;
wire na8246_10;
wire na8248_10;
wire na8250_10;
wire na8252_10;
wire na8254_10;
wire na8256_10;
wire na8258_10;
wire na8262_10;
wire na8263_10;
wire na8264_10;
wire na8266_10;
wire na8269_10;
wire na8273_10;
wire na8279_10;
wire na8282_10;
wire na8290_10;
wire na8293_10;
wire na8299_10;
wire na8303_10;
wire na8308_10;
wire na8316_10;
wire na8321_10;
wire na8331_10;
wire na8335_10;
wire na8340_10;
wire na8350_10;
wire na8353_10;
wire na8364_10;
wire na8368_10;
wire na8374_10;
wire na8380_10;
wire na8423_10;
wire na8424_10;
wire na8425_10;
wire na8426_10;
wire na8427_10;
wire na8428_10;
wire na8429_10;
wire na8430_10;
wire na8431_10;
wire na8432_10;
wire na8433_10;
wire na8434_10;
wire na8435_10;
wire na8436_10;
wire na8437_10;
wire na8438_10;
wire na8439_10;
wire na8440_10;
wire na8441_10;
wire na8442_10;
wire na8443_10;
wire na8444_10;
wire na8445_10;
wire na8446_10;
wire na8447_10;
wire na8448_10;
wire na8449_10;
wire na8450_10;
wire na8451_10;
wire na8452_10;
wire na8453_10;
wire na8454_10;
wire na8455_10;
wire na8456_10;
wire na8457_10;
wire na8458_10;
wire na8459_10;
wire na8460_10;
wire na8461_10;
wire na8462_10;
wire na8463_10;
wire na8464_10;
wire na8465_10;
wire na8466_10;
wire na8467_10;
wire na8468_10;
wire na8469_10;
wire na8470_10;
wire na8471_10;
wire na8472_10;
wire na8473_10;
wire na8474_10;
wire na8475_10;
wire na8476_10;
wire na8477_10;
wire na8478_10;
wire na8479_10;
wire na8480_10;
wire na8481_10;
wire na8482_10;
wire na8483_10;
wire na8484_10;
wire na8485_10;
wire na8486_10;
wire na8487_10;
wire na8488_10;
wire na8489_10;
wire na8490_10;
wire na8491_10;
wire na8492_10;
wire na8493_10;
wire na8494_10;
wire na8495_10;
wire na8496_10;
wire na8497_10;
wire na8499_10;
wire na8501_10;
wire na8503_10;
wire na8505_10;
wire na8507_10;
wire na8509_10;
wire na8511_10;
wire na8513_10;
wire na8515_10;
wire na8517_10;
wire na8519_10;
wire na8521_10;
wire na8523_10;
wire na8525_10;
wire na8527_10;
wire na8529_10;
wire na8531_10;
wire na8533_10;
wire na8535_10;
wire na8537_10;
wire na8539_10;
wire na8543_10;
wire na8544_10;
wire na8545_10;
wire na8547_10;
wire na8549_10;
wire na8551_10;
wire na8553_10;
wire na8555_10;
wire na8557_10;
wire na8559_10;
wire na8561_10;
wire na8563_10;
wire na8565_10;
wire na8567_10;
wire na8569_10;
wire na8571_10;
wire na8573_10;
wire na8575_10;
wire na8579_10;
wire na8581_10;
wire na8585_10;
wire na8587_10;
wire na8589_10;
wire na8591_10;
wire na8593_10;
wire na8595_10;
wire na8597_10;
wire na8599_10;
wire na8601_10;
wire na8603_10;
wire na8605_10;
wire na8607_10;
wire na8609_10;
wire na8611_10;
wire na8613_10;
wire na8615_10;
wire na8617_10;
wire na8619_10;
wire na8621_10;
wire na8623_10;
wire na8625_10;
wire na8627_10;
wire na8629_10;
wire na8631_10;
wire na8633_10;
wire na8635_10;
wire na8637_10;
wire na8639_10;
wire na8641_10;
wire na8643_10;
wire na8645_10;
wire na8647_10;
wire na8649_10;
wire na8651_10;
wire na8653_10;
wire na8655_10;
wire na8657_10;
wire na8659_10;
wire na8661_10;
wire na8663_10;
wire na8665_10;
wire na8667_10;
wire na8671_10;
wire na8672_10;
wire na8673_10;
wire na8675_10;
wire na8677_10;
wire na8679_10;
wire na8681_10;
wire na8683_10;
wire na8685_10;
wire na8687_10;
wire na8689_10;
wire na8691_10;
wire na8693_10;
wire na8695_10;
wire na8697_10;
wire na8699_10;
wire na8701_10;
wire na8703_10;
wire na8707_10;
wire na8709_10;
wire na8713_10;
wire na8715_10;
wire na8717_10;
wire na8719_10;
wire na8721_10;
wire na8723_10;
wire na8725_10;
wire na8727_10;
wire na8729_10;
wire na8731_10;
wire na8733_10;
wire na8735_10;
wire na8737_10;
wire na8739_10;
wire na8741_10;
wire na8743_10;
wire na8745_10;
wire na8747_10;
wire na8749_10;
wire na8751_10;
wire na8753_10;
wire na8755_10;
wire na8757_10;
wire na8759_10;
wire na8761_10;
wire na8763_10;
wire na8765_10;
wire na8767_10;
wire na8769_10;
wire na8771_10;
wire na8773_10;
wire na8775_10;
wire na8777_10;
wire na8779_10;
wire na8781_10;
wire na8783_10;
wire na8785_10;
wire na8787_10;
wire na8789_10;
wire na8791_10;
wire na8793_10;
wire na8795_10;
wire na8798_10;
wire na8799_10;
wire na8801_10;
wire na8803_10;
wire na8805_10;
wire na8807_10;
wire na8809_10;
wire na8811_10;
wire na8813_10;
wire na8817_10;
wire na8819_10;
wire na8821_10;
wire na8823_10;
wire na8825_10;
wire na8827_10;
wire na8829_10;
wire na8831_10;
wire na8833_10;
wire na8835_10;
wire na8837_10;
wire na8839_10;
wire na8841_10;
wire na8843_10;
wire na8845_10;
wire na8847_10;
wire na8849_10;
wire na8851_10;
wire na8853_10;
wire na8855_10;
wire na8857_10;
wire na8859_10;
wire na8863_10;
wire na8864_10;
wire na8865_10;
wire na8867_10;
wire na8869_10;
wire na8871_10;
wire na8873_10;
wire na8875_10;
wire na8877_10;
wire na8879_10;
wire na8881_10;
wire na8883_10;
wire na8885_10;
wire na8887_10;
wire na8889_10;
wire na8891_10;
wire na8893_10;
wire na8895_10;
wire na8899_10;
wire na8901_10;
wire na8905_10;
wire na8907_10;
wire na8909_10;
wire na8911_10;
wire na8913_10;
wire na8915_10;
wire na8917_10;
wire na8919_10;
wire na8921_10;
wire na8923_10;
wire na8925_10;
wire na8927_10;
wire na8929_10;
wire na8931_10;
wire na8933_10;
wire na8935_10;
wire na8937_10;
wire na8939_10;
wire na8941_10;
wire na8943_10;
wire na8945_10;
wire na8947_10;
wire na8949_10;
wire na8951_10;
wire na8953_10;
wire na8955_10;
wire na8957_10;
wire na8959_10;
wire na8961_10;
wire na8963_10;
wire na8965_10;
wire na8967_10;
wire na8969_10;
wire na8971_10;
wire na8973_10;
wire na8975_10;
wire na8977_10;
wire na8979_10;
wire na8981_10;
wire na8983_10;
wire na8985_10;
wire na8987_10;
wire na8991_10;
wire na8992_10;
wire na8993_10;
wire na8995_10;
wire na8997_10;
wire na8999_10;
wire na9001_10;
wire na9003_10;
wire na9005_10;
wire na9007_10;
wire na9009_10;
wire na9011_10;
wire na9013_10;
wire na9015_10;
wire na9017_10;
wire na9019_10;
wire na9021_10;
wire na9023_10;
wire na9025_10;
wire na9027_10;
wire na9029_10;
wire na9031_10;
wire na9033_10;
wire na9035_10;
wire na9037_10;
wire na9039_10;
wire na9041_10;
wire na9043_10;
wire na9045_10;
wire na9047_10;
wire na9049_10;
wire na9051_10;
wire na9053_10;
wire na9055_10;
wire na9057_10;
wire na9059_10;
wire na9061_10;
wire na9063_10;
wire na9065_10;
wire na9067_10;
wire na9069_10;
wire na9071_10;
wire na9073_10;
wire na9075_10;
wire na9077_10;
wire na9079_10;
wire na9081_10;
wire na9083_10;
wire na9085_10;
wire na9087_10;
wire na9089_10;
wire na9091_10;
wire na9093_10;
wire na9095_10;
wire na9097_10;
wire na9099_10;
wire na9101_10;
wire na9103_10;
wire na9105_10;
wire na9107_10;
wire na9109_10;
wire na9111_10;
wire na9113_10;
wire na9115_10;
wire creset_ice40;
wire na6629_109;
wire na6629_110;
wire na6629_111;
wire na6629_112;
wire na6629_113;
wire na6629_114;
wire na6629_115;
wire na6629_116;
wire na6629_117;
wire na6629_118;
wire na6629_119;
wire na6629_120;
wire na6630_100;
wire na6659_100;
wire na6659_113;
wire na6659_114;
wire na6659_115;
wire na6659_116;
wire na6659_117;
wire na6659_118;
wire na6659_119;
wire na6659_120;
wire osc_en_ice40;
wire vio_en_ice40;
wire core_en_ice40;
wire spi_ice40_clk;
wire uart_ice40_rx;
wire uart_ice40_tx;
wire usb_uart_rx;
wire usb_uart_tx;
wire user_led_n0;
wire user_led_n1;
wire user_led_n2;
wire user_led_n3;
wire ice40_io_vio_0;
wire ice40_io_vio_1;
wire ice40_io_vio_2;
wire ice40_io_vio_3;
wire ice40_io_vio_4;
wire ice40_io_vio_5;
wire spi_ice40_cs_n;
wire spi_ice40_miso;
wire spi_ice40_mosi;
wire hyperram_cs_n;
wire hyperram_rwds;
wire spi_flash_clk;
wire hyperram_clk_n;
wire hyperram_clk_p;
wire hyperram_rst_n;
wire ice40_io_vcore_0;
wire ice40_io_vcore_1;
wire ice40_io_vcore_2;
wire ice40_io_vcore_4;
wire spi_flash_cs_n;
wire spi_flash_miso;
wire spi_flash_mosi;
wire power_fauld_ice40;
wire uart_logging_rx;
wire uart_logging_tx;
wire gatemate_debug_3;
wire gatemate_debug_4;
wire gatemate_debug_5;

// C_AND////      x104y101     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1870_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6626_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y56     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2833_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6626_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y102     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3_1 ( .OUT(na3_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1870_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6626_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y55     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4_4 ( .OUT(na4_2), .IN1(na2833_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y49     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na425_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na455_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y50     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6_4 ( .OUT(na6_2), .IN1(na2697_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2695_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x100y81     80'h00_0078_00_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9_1), .IN6(na31_2), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8_4 ( .OUT(na8_2), .IN1(1'b1), .IN2(na450_2), .IN3(na430_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y71     80'h00_0018_00_0000_0888_C888
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9_1 ( .OUT(na9_1), .IN1(na26_2), .IN2(na12_1), .IN3(na469_2), .IN4(na21_1), .IN5(na19_1), .IN6(na13_1), .IN7(1'b1), .IN8(na20_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x85y78     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1502_2), .IN4(~na2439_2), .IN5(1'b1), .IN6(na2773_1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y80     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9675_2), .IN5(~na2440_2), .IN6(1'b0), .IN7(~na807_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x79y76     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1), .IN1(~na811_2), .IN2(~na9610_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2773_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x82y76     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na9675_2), .IN5(~na819_2), .IN6(1'b0), .IN7(~na2442_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y79     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2443_2), .IN8(~na815_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y76     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2444_2), .IN8(~na823_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y77     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na799_2), .IN6(~na2437_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x82y78     80'h00_0018_00_0040_0C33_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1), .IN1(~na803_2), .IN2(~na2438_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2773_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x84y78     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a21_1 ( .OUT(na21_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9139_2), .IN6(na24_1), .IN7(na22_1), .IN8(na23_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x80y81     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na828_2), .IN4(~na2446_2), .IN5(1'b1), .IN6(na2773_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y76     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9341_2), .IN8(~na2447_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y76     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2445_2), .IN8(~na9515_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x83y84     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2448_2), .IN4(~na1494_2), .IN5(1'b1), .IN6(~na2773_1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y75     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a26_4 ( .OUT(na26_2), .IN1(~na29_1), .IN2(~na27_1), .IN3(~na30_1), .IN4(~na28_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y74     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2449_2), .IN8(~na9342_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y78     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9346_2), .IN8(~na2450_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y79     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a29_1 ( .OUT(na29_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2451_2), .IN6(~na9343_2), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x82y81     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2390_2), .IN8(~na863_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y74     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a31_4 ( .OUT(na31_2), .IN1(~na32_1), .IN2(1'b1), .IN3(~na1113_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y73     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na712_1), .IN6(na2773_1), .IN7(~na34_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x80y71     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a34_4 ( .OUT(na34_2), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b1), .IN4(na523_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x75y64     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1), .IN1(na749_2), .IN2(na9605_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2773_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y72     80'h00_0078_00_0000_0C88_C8A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9_1), .IN6(na31_2), .IN7(1'b1), .IN8(na37_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a36_4 ( .OUT(na36_2), .IN1(na9_1), .IN2(na31_2), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y64     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9327_2), .IN8(na2426_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x78y66     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na9675_2), .IN5(na1552_2), .IN6(1'b0), .IN7(na2428_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x90y68     80'h00_0018_00_0000_0888_FCEA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1), .IN1(na9_1), .IN2(1'b0), .IN3(na9144_2), .IN4(na39_1), .IN5(1'b0), .IN6(na31_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x66y74     80'h00_0060_00_0000_0C0E_FFCC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a42_4 ( .OUT(na42_2), .IN1(1'b0), .IN2(na43_1), .IN3(1'b0), .IN4(na6663_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x67y76     80'h00_F618_00_0000_0888_ACFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1), .IN1(na353_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5977_1), .IN7(na517_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a43_5 ( .OUT(na43_2), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na43_1) );
// C_ORAND////      x69y74     80'h00_0018_00_0000_0C88_D3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na43_1), .IN7(~na47_2), .IN8(na42_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x67y80     80'h00_F600_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na47_2), .IN8(~na42_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a46_2 ( .OUT(na46_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na46_1_i) );
// C_///AND/      x70y85     80'h00_0060_00_0000_0C08_FF2C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a47_4 ( .OUT(na47_2), .IN1(1'b1), .IN2(na9246_2), .IN3(na3321_1), .IN4(~na3323_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x64y76     80'h00_0018_00_0000_0888_FEAA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1), .IN1(na6664_1), .IN2(1'b0), .IN3(na517_1), .IN4(1'b0), .IN5(na3328_1), .IN6(na3270_1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x57y71     80'h00_0078_00_0000_0C88_F88F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na51_1), .IN6(na6666_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a50_4 ( .OUT(na50_2), .IN1(1'b1), .IN2(1'b1), .IN3(na53_1), .IN4(na6668_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y71     80'h00_0018_00_0040_0ACF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na5228_2), .IN8(~na5961_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y77     80'h00_0018_00_0040_0ACF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na9865_2), .IN8(~na5962_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y78     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na48_1), .IN5(na3328_1), .IN6(1'b0), .IN7(na6671_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y102     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a56_4 ( .OUT(na56_2), .IN1(na971_1), .IN2(~na1358_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y52     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1223_1), .IN8(na973_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x105y52     80'h00_FA00_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1_i), .IN1(na6672_1), .IN2(1'b0), .IN3(na1223_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na973_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_2 ( .OUT(na58_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na58_1_i) );
// C_MX2b////      x99y52     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na973_1), .IN5(na2991_1), .IN6(1'b0), .IN7(na1223_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y60     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2423_2), .IN8(na9323_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y61     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(na741_2), .IN6(na9604_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x99y70     80'h00_0018_00_0040_0AB3_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1), .IN1(1'b1), .IN2(~na36_2), .IN3(1'b1), .IN4(na6673_2), .IN5(~na9944_2), .IN6(~na36_1), .IN7(1'b0),
                    .IN8(na6674_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x78y65     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2424_2), .IN4(na9326_2), .IN5(1'b1), .IN6(~na2773_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x93y76     80'h00_0078_00_0000_0C88_D5CD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9947_2), .IN6(1'b0), .IN7(~na9148_2), .IN8(na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a67_4 ( .OUT(na67_2), .IN1(~na9237_2), .IN2(na36_1), .IN3(1'b0), .IN4(na41_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y69     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a68_4 ( .OUT(na68_2), .IN1(1'b1), .IN2(na36_2), .IN3(1'b1), .IN4(~na6673_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x91y72     80'h00_0018_00_0040_0C26_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1), .IN1(1'b0), .IN2(~na9946_2), .IN3(na6675_2), .IN4(1'b0), .IN5(1'b1), .IN6(na36_1), .IN7(1'b1), .IN8(na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x100y68     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9947_2), .IN6(1'b0), .IN7(~na9148_2), .IN8(~na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x100y69     80'h00_0018_00_0040_0C15_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a71_1 ( .OUT(na71_1), .IN1(~na9947_2), .IN2(1'b0), .IN3(na9148_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y67     80'h00_0018_00_0040_0AB5_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_1 ( .OUT(na72_1), .IN1(1'b1), .IN2(~na36_2), .IN3(1'b1), .IN4(na6673_2), .IN5(~na9947_2), .IN6(na6677_2), .IN7(1'b1),
                    .IN8(na6678_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y68     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na36_2), .IN7(1'b1), .IN8(na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x103y66     80'h00_0018_00_0040_0AF6_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1), .IN1(1'b1), .IN2(~na36_2), .IN3(1'b1), .IN4(na6673_2), .IN5(na9947_2), .IN6(~na36_1), .IN7(~na9145_2),
                    .IN8(na6674_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y68     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9947_2), .IN6(1'b1), .IN7(1'b1), .IN8(na73_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x100y65     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a76_4 ( .OUT(na76_2), .IN1(1'b0), .IN2(na36_2), .IN3(1'b0), .IN4(~na6673_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x99y67     80'h00_0060_00_0000_0C08_FFC9
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a77_4 ( .OUT(na77_2), .IN1(na9947_2), .IN2(na36_2), .IN3(1'b0), .IN4(~na6673_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x101y64     80'h00_0018_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9947_2), .IN6(na36_2), .IN7(1'b0), .IN8(~na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x100y73     80'h00_0018_00_0040_0C26_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1), .IN1(1'b0), .IN2(~na6681_1), .IN3(na6675_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na36_1), .IN7(1'b1), .IN8(na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x102y74     80'h00_0018_00_0040_0C4E_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1), .IN1(1'b0), .IN2(na36_1), .IN3(~na6684_1), .IN4(na6673_2), .IN5(na9947_2), .IN6(1'b1), .IN7(1'b1),
                    .IN8(na9149_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x94y69     80'h00_0078_00_0000_0C88_A5AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9947_2), .IN6(1'b1), .IN7(na82_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a81_4 ( .OUT(na81_2), .IN1(1'b1), .IN2(na35_1), .IN3(na8_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y65     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a82_1 ( .OUT(na82_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na36_2), .IN7(1'b1), .IN8(~na6673_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x104y73     80'h00_FE00_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na478_2), .IN8(na6466_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a83_2 ( .OUT(na83_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na83_1_i) );
// C_MX2b////      x76y63     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(na9606_2), .IN6(na759_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y60     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2430_2), .IN6(na763_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x79y67     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1), .IN1(na2431_2), .IN2(na9331_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2773_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y70     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2432_2), .IN6(na9332_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x75y63     80'h00_FE18_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(na9607_2), .IN6(na9333_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a88_5 ( .OUT(na88_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na88_1) );
// C_MX2b////D      x71y66     80'h00_FE18_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9608_2), .IN8(na779_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a89_5 ( .OUT(na89_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1) );
// C_MX2b////D      x80y65     80'h00_FE18_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2435_2), .IN6(na786_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_5 ( .OUT(na90_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1) );
// C_MX2a////D      x81y58     80'h00_FE18_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a91_1 ( .OUT(na91_1), .IN1(na2436_2), .IN2(na792_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2773_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a91_5 ( .OUT(na91_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na91_1) );
// C_AND///AND/      x102y86     80'h00_0078_00_0000_0C88_3C48
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2768_2), .IN7(1'b1), .IN8(~na2820_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a92_4 ( .OUT(na92_2), .IN1(na2960_1), .IN2(na758_2), .IN3(~na757_1), .IN4(na783_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x93y81     80'h00_0078_00_0000_0C88_4525
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a95_1 ( .OUT(na95_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2960_1), .IN6(1'b1), .IN7(~na757_1), .IN8(na783_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a95_4 ( .OUT(na95_2), .IN1(~na2960_1), .IN2(1'b1), .IN3(na757_1), .IN4(~na783_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x88y83     80'h00_0078_00_0000_0C88_8515
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2960_1), .IN6(1'b1), .IN7(na757_1), .IN8(na783_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a97_4 ( .OUT(na97_2), .IN1(~na2960_1), .IN2(1'b1), .IN3(~na757_1), .IN4(~na783_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x101y88     80'h00_0060_00_0000_0C06_FFC3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a99_4 ( .OUT(na99_2), .IN1(1'b0), .IN2(~na2768_2), .IN3(1'b0), .IN4(na2820_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x95y89     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a100_4 ( .OUT(na100_2), .IN1(~na95_2), .IN2(~na2780_1), .IN3(~na2740_1), .IN4(~na101_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x88y86     80'h00_0060_00_0000_0C08_FFEA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a101_4 ( .OUT(na101_2), .IN1(na2960_1), .IN2(1'b0), .IN3(na757_1), .IN4(na783_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y83     80'h00_0018_00_0000_0C88_1CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2894_2), .IN7(~na2838_1), .IN8(~na2836_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x109y91     80'h00_FA18_00_0000_0888_4FFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1), .IN1(1'b1), .IN2(na2894_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2838_1), .IN8(na2836_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a103_5 ( .OUT(na103_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na103_1) );
// C_MX4b////      x91y70     80'h00_0018_00_0040_0A3F_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1), .IN1(1'b1), .IN2(na2935_1), .IN3(na2937_2), .IN4(1'b1), .IN5(~na919_1), .IN6(~na1083_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y89     80'h00_0078_00_0000_0C88_2CAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2894_2), .IN7(na2838_1), .IN8(~na2836_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a106_4 ( .OUT(na106_2), .IN1(1'b1), .IN2(na99_2), .IN3(na102_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x106y90     80'h00_FA18_00_0000_0788_7F7D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a107_1 ( .OUT(na107_1), .IN1(~na103_1), .IN2(na6695_1), .IN3(~na106_1), .IN4(~na6468_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na106_2),
                     .IN8(~na6696_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a107_5 ( .OUT(na107_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na107_1) );
// C_///AND/      x87y79     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a112_4 ( .OUT(na112_2), .IN1(na95_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na16_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y76     80'h00_0018_00_0040_0A3F_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a114_1 ( .OUT(na114_1), .IN1(1'b1), .IN2(na2935_1), .IN3(na2937_2), .IN4(1'b1), .IN5(~na918_1), .IN6(~na1082_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x110y90     80'h00_FA18_00_0000_0788_7F7D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a116_1 ( .OUT(na116_1), .IN1(~na103_1), .IN2(na6705_1), .IN3(~na106_1), .IN4(~na6469_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na106_2),
                     .IN8(~na6706_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a116_5 ( .OUT(na116_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na116_1) );
// C_///AND/      x84y78     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a120_4 ( .OUT(na120_2), .IN1(~na17_1), .IN2(1'b1), .IN3(na9170_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x91y81     80'h00_0018_00_0040_0A3F_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(1'b1), .IN2(na2935_1), .IN3(na2937_2), .IN4(1'b1), .IN5(~na917_1), .IN6(~na9395_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x78y72     80'h00_0018_00_0000_0888_D77D
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1), .IN1(~na95_1), .IN2(na18_1), .IN3(~na97_1), .IN4(~na39_1), .IN5(~na95_2), .IN6(~na91_1), .IN7(~na97_2),
                     .IN8(na9142_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x94y81     80'h00_0018_00_0040_0AAF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(na2937_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na916_1), .IN7(1'b1),
                     .IN8(~na963_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x105y87     80'h00_FA18_00_0000_0788_FD7D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a129_1 ( .OUT(na129_1), .IN1(~na9178_2), .IN2(na6719_1), .IN3(~na106_1), .IN4(~na6471_1), .IN5(~na103_1), .IN6(na6723_1),
                     .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a129_5 ( .OUT(na129_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na129_1) );
// C_MX4b////      x89y81     80'h00_0018_00_0040_0ACF_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(~na2937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2970_1),
                     .IN8(~na9351_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x110y89     80'h00_FA18_00_0000_0788_DF7D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a135_1 ( .OUT(na135_1), .IN1(~na103_1), .IN2(na9949_2), .IN3(~na106_1), .IN4(~na6472_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na102_1),
                     .IN8(na6727_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a135_5 ( .OUT(na135_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na135_1) );
// C_ORAND////      x81y81     80'h00_0018_00_0000_0888_FDD7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(~na9173_2), .IN2(~na85_1), .IN3(~na9172_2), .IN4(na20_1), .IN5(~na95_1), .IN6(na9138_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y85     80'h00_0018_00_0040_0ACF_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(~na2937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1005_1),
                     .IN8(~na2967_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x109y90     80'h00_FA18_00_0000_0788_F37D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(~na103_1), .IN2(na6736_2), .IN3(~na106_1), .IN4(~na6473_1), .IN5(1'b0), .IN6(~na144_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a142_5 ( .OUT(na142_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na142_1) );
// C_ORAND////      x101y84     80'h00_0018_00_0000_0888_FEA5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a144_1 ( .OUT(na144_1), .IN1(~na145_1), .IN2(1'b0), .IN3(na102_1), .IN4(1'b0), .IN5(na9176_2), .IN6(na99_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x93y83     80'h00_0018_00_0000_0888_D7DC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a145_1 ( .OUT(na145_1), .IN1(1'b0), .IN2(na99_2), .IN3(~na9170_2), .IN4(na23_1), .IN5(~na86_1), .IN6(~na9174_2), .IN7(~na9172_2),
                     .IN8(na9135_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x93y82     80'h00_0018_00_0040_0ACF_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a147_1 ( .OUT(na147_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(~na2937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1004_1),
                     .IN8(~na838_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x108y91     80'h00_FA18_00_0000_0788_FD7C
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a149_1 ( .OUT(na149_1), .IN1(1'b0), .IN2(na6743_1), .IN3(~na106_1), .IN4(~na6474_1), .IN5(~na103_1), .IN6(na6749_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a149_5 ( .OUT(na149_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na149_1) );
// C_MX4b////      x97y75     80'h00_0018_00_0040_0A92_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a151_1 ( .OUT(na151_1), .IN1(~na9176_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na152_1), .IN5(na6745_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(na154_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y82     80'h00_0018_00_0000_0888_FD7D
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(~na95_2), .IN2(na13_1), .IN3(~na97_1), .IN4(~na87_1), .IN5(~na95_1), .IN6(na25_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x104y80     80'h00_0078_00_0000_0C88_C3C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2768_2), .IN7(1'b1), .IN8(na2820_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a154_4 ( .OUT(na154_2), .IN1(~na2981_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6752_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y75     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2773_1), .IN7(1'b1), .IN8(na5585_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y104     80'h00_0018_00_0040_0ACF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(1'b1), .IN2(na2935_1), .IN3(~na2937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2966_1),
                     .IN8(~na1003_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x98y82     80'h00_FE18_00_0000_0888_5FFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a159_1 ( .OUT(na159_1), .IN1(1'b1), .IN2(na5586_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a159_5 ( .OUT(na159_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na159_1) );
// C_MX4b/D///      x104y76     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_1 ( .OUT(na160_1_i), .IN1(1'b1), .IN2(na161_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9181_2), .IN6(na6479_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_2 ( .OUT(na160_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na160_1_i) );
// C_///AND/      x101y76     80'h00_0060_00_0000_0C08_FF2A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a161_4 ( .OUT(na161_2), .IN1(na8107_2), .IN2(1'b1), .IN3(na2950_1), .IN4(~na2948_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x103y74     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1_i), .IN1(1'b1), .IN2(~na161_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na6480_1), .IN6(na164_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_2 ( .OUT(na164_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na164_1_i) );
// C_MX4b/D///      x102y78     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_1 ( .OUT(na165_1_i), .IN1(1'b1), .IN2(na161_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9182_2), .IN6(na6481_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_2 ( .OUT(na165_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na165_1_i) );
// C_MX4b/D///      x106y80     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1_i), .IN1(1'b1), .IN2(na161_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9183_2), .IN6(na6482_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_2 ( .OUT(na166_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na166_1_i) );
// C_MX4b/D///      x107y78     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_1 ( .OUT(na167_1_i), .IN1(1'b1), .IN2(~na161_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na6484_1), .IN6(na167_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_2 ( .OUT(na167_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na167_1_i) );
// C_MX4b/D///      x103y79     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1_i), .IN1(1'b1), .IN2(na169_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na168_1), .IN6(na6477_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_2 ( .OUT(na168_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na168_1_i) );
// C_///AND/      x107y80     80'h00_0060_00_0000_0C08_FF4A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a169_4 ( .OUT(na169_2), .IN1(na8107_2), .IN2(1'b1), .IN3(~na2950_1), .IN4(na2948_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x102y77     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_1 ( .OUT(na170_1_i), .IN1(1'b1), .IN2(na169_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na170_1),
                     .IN8(na6478_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_2 ( .OUT(na170_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na170_1_i) );
// C_AND*/D///      x91y50     80'h00_FE00_00_0000_0388_3CFF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a171_1 ( .OUT(na171_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(1'b1), .IN8(~na4091_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a171_2 ( .OUT(na171_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na171_1_i) );
// C_///AND/      x91y54     80'h00_0060_00_0000_0C08_FF34
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a172_4 ( .OUT(na172_2), .IN1(~na32_1), .IN2(na173_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y78     80'h00_0018_00_0000_0888_134F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1113_2), .IN4(na174_1), .IN5(1'b1), .IN6(~na2252_1), .IN7(~na1113_1),
                     .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x98y78     80'h00_0018_00_0000_0888_FD55
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a174_1 ( .OUT(na174_1), .IN1(~na214_1), .IN2(1'b0), .IN3(~na210_1), .IN4(1'b0), .IN5(~na214_2), .IN6(na9179_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x86y60     80'h00_0018_00_0000_0888_9999
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(~na88_1), .IN2(~na3731_2), .IN3(~na9852_2), .IN4(~na87_1), .IN5(na3703_2), .IN6(na9165_2), .IN7(na84_1),
                     .IN8(na9850_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x88y66     80'h00_0060_00_0000_0C06_FF5C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a178_4 ( .OUT(na178_2), .IN1(1'b0), .IN2(na3727_2), .IN3(~na84_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x83y66     80'h00_0018_00_0000_0C66_5A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3703_2), .IN6(1'b0), .IN7(~na90_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x88y65     80'h00_0078_00_0000_0C66_3306
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3731_1), .IN7(1'b0), .IN8(~na87_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a180_4 ( .OUT(na180_2), .IN1(~na88_1), .IN2(~na3731_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x89y66     80'h00_0018_00_0000_0888_9956
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(na3707_1), .IN2(~na6759_1), .IN3(na9846_2), .IN4(1'b0), .IN5(na3729_1), .IN6(na85_1), .IN7(na9835_2),
                     .IN8(na9162_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x87y63     80'h00_0018_00_0000_0888_9F69
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(~na3725_1), .IN2(~na9150_2), .IN3(na420_1), .IN4(~na61_1), .IN5(1'b0), .IN6(1'b0), .IN7(na66_1),
                     .IN8(na9842_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x87y61     80'h00_0018_00_0000_0888_9A99
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a189_1 ( .OUT(na189_1), .IN1(~na3725_2), .IN2(~na35_1), .IN3(~na63_1), .IN4(~na9843_2), .IN5(~na193_1), .IN6(1'b0), .IN7(na9849_2),
                     .IN8(na39_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y67     80'h00_0018_00_0040_0A32_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(na9853_2), .IN5(na6767_2), .IN6(~na2962_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y74     80'h00_0018_00_0000_0888_8438
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(na29_1), .IN2(na27_1), .IN3(1'b1), .IN4(~na28_1), .IN5(~na32_1), .IN6(na18_1), .IN7(na30_1),
                     .IN8(na21_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y65     80'h00_0018_00_0000_0888_1283
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a197_1 ( .OUT(na197_1), .IN1(1'b1), .IN2(~na3714_1), .IN3(na199_1), .IN4(na207_1), .IN5(na203_1), .IN6(~na3718_1), .IN7(~na9845_2),
                     .IN8(~na9848_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x94y67     80'h00_0018_00_0000_0888_6663
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1), .IN1(1'b0), .IN2(na3722_1), .IN3(~na6769_1), .IN4(na9838_2), .IN5(~na6770_1), .IN6(na3705_2), .IN7(na9837_2),
                     .IN8(~na6768_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x91y63     80'h00_0018_00_0000_0888_6939
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a203_1 ( .OUT(na203_1), .IN1(na86_1), .IN2(na9851_2), .IN3(1'b0), .IN4(na9847_2), .IN5(na9836_2), .IN6(na91_1), .IN7(na9841_2),
                     .IN8(~na6771_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x94y70     80'h00_0018_00_0000_0888_6A65
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(na3716_1), .IN2(1'b0), .IN3(na9840_2), .IN4(~na6775_1), .IN5(~na3720_1), .IN6(1'b0), .IN7(~na6774_1),
                     .IN8(na9839_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y73     80'h00_0018_00_0000_0888_C888
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a210_1 ( .OUT(na210_1), .IN1(na186_1), .IN2(na211_2), .IN3(na197_1), .IN4(na194_1), .IN5(na189_1), .IN6(na182_1), .IN7(1'b1),
                     .IN8(na177_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y86     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a211_4 ( .OUT(na211_2), .IN1(na212_1), .IN2(na2935_1), .IN3(na2937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y87     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7054_2), .IN6(1'b1), .IN7(na9177_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y73     80'h00_0078_00_0000_0C88_3882
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na155_1), .IN6(na215_1), .IN7(1'b1), .IN8(~na154_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a214_4 ( .OUT(na214_2), .IN1(na2920_2), .IN2(~na2894_2), .IN3(na2838_1), .IN4(na2836_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y90     80'h00_0018_00_0000_0888_8282
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a215_1 ( .OUT(na215_1), .IN1(na223_1), .IN2(~na6778_1), .IN3(na220_1), .IN4(na753_2), .IN5(na6776_1), .IN6(~na6778_2), .IN7(na6777_2),
                     .IN8(na6779_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y99     80'h00_0018_00_0000_0888_53A2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1), .IN1(na6783_1), .IN2(~na6782_2), .IN3(na6780_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na6781_1), .IN7(~na6784_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y89     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a223_1 ( .OUT(na223_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7054_2), .IN6(1'b1), .IN7(na224_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y89     80'h00_0018_00_0000_0C88_23FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2894_2), .IN7(na2838_1), .IN8(~na2836_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y64     80'h00_0018_00_0000_0888_2128
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a228_1 ( .OUT(na228_1), .IN1(na234_2), .IN2(na233_1), .IN3(na232_1), .IN4(~na2901_1), .IN5(~na2902_1), .IN6(~na2904_1), .IN7(na232_2),
                     .IN8(~na2901_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y53     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2900_2), .IN6(~na2898_2), .IN7(~na2899_2),
                     .IN8(~na2897_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a232_4 ( .OUT(na232_2), .IN1(~na2900_1), .IN2(~na2898_1), .IN3(~na2899_1), .IN4(~na2897_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y52     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na281_2), .IN6(~na171_1), .IN7(~na300_1), .IN8(~na301_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y51     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a234_4 ( .OUT(na234_2), .IN1(~na2917_2), .IN2(~na2904_2), .IN3(~na9705_2), .IN4(~na2907_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x101y71     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_1 ( .OUT(na235_1_i), .IN1(1'b1), .IN2(na169_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na235_1), .IN6(na6479_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_2 ( .OUT(na235_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na235_1_i) );
// C_AND////D      x112y74     80'h00_FA18_00_0000_0888_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_1 ( .OUT(na236_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4856_1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a236_5 ( .OUT(na236_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na236_1) );
// C_ICOMP////      x114y78     80'h00_0018_00_0000_0888_3FC6
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(~na4894_1), .IN2(na9864_2), .IN3(1'b0), .IN4(~na6476_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na238_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x116y96     80'h00_0060_00_0000_0C08_FF51
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a238_4 ( .OUT(na238_2), .IN1(~na995_1), .IN2(~na2671_1), .IN3(~na2673_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x111y74     80'h00_FA18_00_0000_0888_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(1'b1), .IN2(na4861_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a239_5 ( .OUT(na239_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na239_1) );
// C_AND////D      x111y76     80'h00_FA18_00_0000_0888_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_1 ( .OUT(na240_1), .IN1(1'b1), .IN2(1'b1), .IN3(na4865_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a240_5 ( .OUT(na240_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na240_1) );
// C_AND////D      x111y75     80'h00_FA18_00_0000_0888_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_1 ( .OUT(na241_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4869_1), .IN6(1'b1), .IN7(1'b1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a241_5 ( .OUT(na241_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na241_1) );
// C_AND////D      x113y76     80'h00_FA18_00_0000_0888_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a242_1 ( .OUT(na242_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4873_1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a242_5 ( .OUT(na242_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na242_1) );
// C_AND////D      x109y73     80'h00_FA18_00_0000_0888_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4878_1), .IN7(1'b1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a243_5 ( .OUT(na243_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na243_1) );
// C_AND////D      x110y73     80'h00_FA18_00_0000_0888_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a244_1 ( .OUT(na244_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a244_5 ( .OUT(na244_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na244_1) );
// C_AND////D      x110y75     80'h00_FA18_00_0000_0888_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a245_1 ( .OUT(na245_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4887_1), .IN6(1'b1), .IN7(1'b1), .IN8(na237_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a245_5 ( .OUT(na245_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na245_1) );
// C_MX4b/D///      x101y74     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_1 ( .OUT(na246_1_i), .IN1(1'b1), .IN2(~na169_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na6480_1), .IN6(na246_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_2 ( .OUT(na246_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na246_1_i) );
// C_MX4b/D///      x100y105     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_1 ( .OUT(na247_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na247_1),
                     .IN8(na3757_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_2 ( .OUT(na247_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na247_1_i) );
// C_///AND/      x101y103     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a248_4 ( .OUT(na248_2), .IN1(1'b1), .IN2(1'b1), .IN3(na9188_2), .IN4(~na6786_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x99y101     80'h00_0078_00_0000_0C88_8888
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a251_1 ( .OUT(na251_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9764_2), .IN6(na3138_1), .IN7(na3134_1), .IN8(na3139_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a251_4 ( .OUT(na251_2), .IN1(na3169_1), .IN2(na3170_1), .IN3(na3190_1), .IN4(na3192_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y104     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3208_1), .IN6(na3205_1), .IN7(na3195_1), .IN8(na3201_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y104     80'h00_0018_00_0000_0888_888C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(1'b1), .IN2(na256_2), .IN3(na2157_1), .IN4(na257_1), .IN5(na1903_1), .IN6(na258_2), .IN7(na1829_1),
                     .IN8(na2255_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y104     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a256_4 ( .OUT(na256_2), .IN1(na1695_1), .IN2(na1656_1), .IN3(na247_1), .IN4(na322_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y104     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a257_1 ( .OUT(na257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3118_1), .IN6(na3126_1), .IN7(na3113_1), .IN8(na3119_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y104     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a258_4 ( .OUT(na258_2), .IN1(na2721_1), .IN2(na2895_1), .IN3(na2748_1), .IN4(na2739_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x101y80     80'h00_FE18_00_0000_0888_5FCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a259_1 ( .OUT(na259_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a259_5 ( .OUT(na259_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na259_1) );
// C_AND////D      x104y79     80'h00_FE18_00_0000_0888_5FFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1), .IN1(1'b1), .IN2(na5588_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a260_5 ( .OUT(na260_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na260_1) );
// C_AND////D      x104y77     80'h00_FE18_00_0000_0888_5FAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a261_1 ( .OUT(na261_1), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a261_5 ( .OUT(na261_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na261_1) );
// C_AND////D      x99y82     80'h00_FE18_00_0000_0888_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a262_5 ( .OUT(na262_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na262_1) );
// C_AND////D      x100y83     80'h00_FE18_00_0000_0888_5FFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a263_1 ( .OUT(na263_1), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a263_5 ( .OUT(na263_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na263_1) );
// C_AND////D      x102y83     80'h00_FE18_00_0000_0888_5FFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a264_1 ( .OUT(na264_1), .IN1(1'b1), .IN2(na5592_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a264_5 ( .OUT(na264_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na264_1) );
// C_AND////D      x105y82     80'h00_FE18_00_0000_0888_5FFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a265_5 ( .OUT(na265_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na265_1) );
// C_MX4b/D///      x105y71     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_1 ( .OUT(na266_1_i), .IN1(1'b1), .IN2(na169_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na266_1), .IN6(na6481_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_2 ( .OUT(na266_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na266_1_i) );
// C_MX4b/D///      x105y78     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1_i), .IN1(na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9189_2),
                     .IN8(na6478_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_2 ( .OUT(na267_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na267_1_i) );
// C_AND////      x103y73     80'h00_0018_00_0000_0C88_1AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_1 ( .OUT(na268_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8107_2), .IN6(1'b1), .IN7(~na2950_1), .IN8(~na2948_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x97y79     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_1 ( .OUT(na269_1_i), .IN1(1'b1), .IN2(na169_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na269_1), .IN6(na6482_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_2 ( .OUT(na269_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na269_1_i) );
// C_MX4b/D///      x103y77     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a270_1 ( .OUT(na270_1_i), .IN1(1'b1), .IN2(na169_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na270_1), .IN6(na6483_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a270_2 ( .OUT(na270_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na270_1_i) );
// C_MX4b/D///      x103y76     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_1 ( .OUT(na271_1_i), .IN1(1'b1), .IN2(~na169_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na6484_1), .IN6(na271_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_2 ( .OUT(na271_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na271_1_i) );
// C_MX4b/D///      x94y100     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1_i), .IN1(1'b1), .IN2(~na273_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na277_1),
                     .IN8(na272_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a272_2 ( .OUT(na272_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na272_1_i) );
// C_AND////      x93y98     80'h00_0018_00_0000_0888_4152
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1), .IN1(na3354_1), .IN2(~na3424_2), .IN3(~na3276_1), .IN4(1'b1), .IN5(~na3588_1), .IN6(~na3299_2), .IN7(~na3301_1),
                     .IN8(na3216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y105     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na278_1), .IN8(~na272_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y103     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na279_1), .IN6(1'b1), .IN7(na282_1), .IN8(na272_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x91y99     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a279_1 ( .OUT(na279_1_i), .IN1(1'b1), .IN2(na273_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na279_1), .IN6(na280_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a279_2 ( .OUT(na279_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na279_1_i) );
// C_///AND/      x93y108     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a280_4 ( .OUT(na280_2), .IN1(1'b1), .IN2(na3903_1), .IN3(~na278_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x91y51     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a281_4 ( .OUT(na281_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(1'b1), .IN4(na4091_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a281_5 ( .OUT(na281_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na281_2_i) );
// C_MX4b/D///      x94y101     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1_i), .IN1(1'b1), .IN2(na273_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na282_1),
                     .IN8(na283_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a282_2 ( .OUT(na282_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na282_1_i) );
// C_///AND/      x92y106     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a283_4 ( .OUT(na283_2), .IN1(1'b1), .IN2(na3903_2), .IN3(~na278_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y101     80'h00_0018_00_0000_0888_1354
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_1 ( .OUT(na285_1), .IN1(~na3588_1), .IN2(na3299_2), .IN3(~na3276_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3424_2), .IN7(~na3301_1),
                     .IN8(~na3216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y113     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na325_2), .IN5(1'b0), .IN6(~na291_2), .IN7(1'b0), .IN8(~na6787_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x86y116     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a288_4 ( .OUT(na288_2), .IN1(na9192_2), .IN2(na291_1), .IN3(na289_2), .IN4(na9193_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x88y111     80'h00_FE00_80_0000_0C88_F135
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a289_1 ( .OUT(na289_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na285_1), .IN6(~na290_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a289_2 ( .OUT(na289_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na289_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a289_4 ( .OUT(na289_2_i), .IN1(~na285_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na294_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a289_5 ( .OUT(na289_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na289_2_i) );
// C_MX2b////      x87y114     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a290_1 ( .OUT(na290_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na325_2), .IN5(~na6788_2), .IN6(1'b0), .IN7(~na289_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x89y112     80'h00_FE00_80_0000_0C88_3555
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a291_1 ( .OUT(na291_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na285_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na292_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a291_2 ( .OUT(na291_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na291_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a291_4 ( .OUT(na291_2_i), .IN1(~na285_1), .IN2(1'b1), .IN3(~na287_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a291_5 ( .OUT(na291_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na291_2_i) );
// C_MX2b////      x86y114     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a292_1 ( .OUT(na292_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na325_2), .IN5(1'b0), .IN6(~na291_1), .IN7(1'b0), .IN8(~na6789_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y116     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a294_1 ( .OUT(na294_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na325_2), .IN5(~na6790_2), .IN6(1'b0), .IN7(~na289_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x106y82     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_1 ( .OUT(na295_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6792_2), .IN6(na299_2), .IN7(1'b0), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_2 ( .OUT(na295_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na295_1_i) );
// C_ORAND////      x111y85     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a296_1 ( .OUT(na296_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6936_2), .IN6(na9194_2), .IN7(1'b0), .IN8(na154_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x110y83     80'h00_0078_00_0000_0C88_428F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a298_1 ( .OUT(na298_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2918_1), .IN6(~na2894_2), .IN7(~na2838_1),
                     .IN8(na2836_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a298_4 ( .OUT(na298_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2838_1), .IN4(na3540_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x109y74     80'h00_0060_00_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a299_4 ( .OUT(na299_2), .IN1(na2924_1), .IN2(1'b1), .IN3(na298_1), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*/D///      x94y51     80'h00_FE00_00_0000_0388_5CFF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a300_1 ( .OUT(na300_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(~na4089_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a300_2 ( .OUT(na300_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na300_1_i) );
// C_///AND/D      x88y48     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a301_4 ( .OUT(na301_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(na4089_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a301_5 ( .OUT(na301_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na301_2_i) );
// C_AND////      x99y98     80'h00_0018_00_0000_0888_512A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a303_1 ( .OUT(na303_1), .IN1(na3297_2), .IN2(1'b1), .IN3(na3357_1), .IN4(~na3423_1), .IN5(~na3297_1), .IN6(~na3600_1), .IN7(~na3292_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x97y105     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a306_1 ( .OUT(na306_1_i), .IN1(1'b1), .IN2(na303_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na306_1), .IN6(na307_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a306_2 ( .OUT(na306_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na306_1_i) );
// C_///AND/      x97y106     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a307_4 ( .OUT(na307_2), .IN1(~na306_1), .IN2(~na308_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y104     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a308_1 ( .OUT(na308_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na306_1), .IN6(na311_1), .IN7(na309_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x98y105     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1_i), .IN1(1'b1), .IN2(na303_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na309_1),
                     .IN8(na310_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a309_2 ( .OUT(na309_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na309_1_i) );
// C_AND////      x98y112     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a310_1 ( .OUT(na310_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na308_1), .IN7(na3896_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x95y106     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1_i), .IN1(1'b1), .IN2(~na303_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na312_2), .IN6(na311_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a311_2 ( .OUT(na311_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na311_1_i) );
// C_///AND/      x97y111     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a312_4 ( .OUT(na312_2), .IN1(1'b1), .IN2(~na308_1), .IN3(na3896_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x97y97     80'h00_FE00_00_0000_0888_1424
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a313_1 ( .OUT(na313_1_i), .IN1(~na9940_2), .IN2(na5223_2), .IN3(na3357_1), .IN4(~na3423_1), .IN5(~na3297_2), .IN6(na3600_1),
                     .IN7(~na3292_1), .IN8(~na9812_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a313_2 ( .OUT(na313_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na313_1_i) );
// C_AND////      x121y112     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_1 ( .OUT(na316_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9935_2), .IN6(na6794_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x131y118     80'h00_F900_80_0000_0C88_ACF2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_1 ( .OUT(na318_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na316_1), .IN7(na4021_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a318_2 ( .OUT(na318_1), .CLK(~na4116_1), .EN(na3238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na318_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a318_4 ( .OUT(na318_2_i), .IN1(na9196_2), .IN2(~na318_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a318_5 ( .OUT(na318_2), .CLK(~na4116_1), .EN(na3238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na318_2_i) );
// C_AND/D//AND/D      x130y119     80'h00_F900_80_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_1 ( .OUT(na320_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na316_1), .IN7(1'b1), .IN8(na4023_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a320_2 ( .OUT(na320_1), .CLK(~na4116_1), .EN(na3238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na320_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a320_4 ( .OUT(na320_2_i), .IN1(1'b1), .IN2(na316_1), .IN3(na4021_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a320_5 ( .OUT(na320_2), .CLK(~na4116_1), .EN(na3238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na320_2_i) );
// C_///AND/D      x136y122     80'h00_F900_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a321_4 ( .OUT(na321_2_i), .IN1(1'b1), .IN2(na316_1), .IN3(1'b1), .IN4(na4023_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a321_5 ( .OUT(na321_2), .CLK(~na4116_1), .EN(na3238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na321_2_i) );
// C_MX4b/D///      x98y106     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3759_2),
                     .IN8(na322_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_2 ( .OUT(na322_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na322_1_i) );
// C_AND////      x89y111     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9940_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na325_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x94y114     80'h00_FE18_00_0000_0888_3F83
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(1'b1), .IN2(~na326_2), .IN3(na333_1), .IN4(na1859_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1859_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a325_5 ( .OUT(na325_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na325_1) );
// C_///AND/D      x87y118     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a326_4 ( .OUT(na326_2_i), .IN1(na324_1), .IN2(na3892_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a326_5 ( .OUT(na326_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na326_2_i) );
// C_AND////      x99y105     80'h00_0018_00_0000_0888_35A1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1), .IN1(~na3297_2), .IN2(~na3600_1), .IN3(na3292_1), .IN4(1'b1), .IN5(~na3297_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na3423_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y114     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a331_1 ( .OUT(na331_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na325_2), .IN5(~na6796_2), .IN6(1'b0), .IN7(~na336_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y113     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a332_4 ( .OUT(na332_2), .IN1(na338_2), .IN2(na334_1), .IN3(na336_1), .IN4(na9200_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x88y119     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a333_1 ( .OUT(na333_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3894_1), .IN6(1'b1), .IN7(1'b1), .IN8(na9199_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a333_2 ( .OUT(na333_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na333_1_i) );
// C_AND/D///      x93y112     80'h00_FE00_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a334_1 ( .OUT(na334_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na329_1), .IN6(1'b1), .IN7(~na335_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a334_2 ( .OUT(na334_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na334_1_i) );
// C_MX2b////      x92y113     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na325_2), .IN5(1'b0), .IN6(~na334_1), .IN7(1'b0), .IN8(~na6797_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x94y111     80'h00_FE00_80_0000_0C88_F135
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a336_1 ( .OUT(na336_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na329_1), .IN6(~na337_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a336_2 ( .OUT(na336_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na336_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a336_4 ( .OUT(na336_2_i), .IN1(~na329_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na331_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a336_5 ( .OUT(na336_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na336_2_i) );
// C_MX2b////      x93y116     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a337_1 ( .OUT(na337_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na325_2), .IN5(~na6798_2), .IN6(1'b0), .IN7(~na336_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x93y113     80'h00_FE00_80_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a338_4 ( .OUT(na338_2_i), .IN1(~na329_1), .IN2(1'b1), .IN3(~na339_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a338_5 ( .OUT(na338_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na338_2_i) );
// C_MX2b////      x90y115     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a339_1 ( .OUT(na339_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na325_2), .IN5(~na338_2), .IN6(1'b0), .IN7(~na6799_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y70     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a340_1 ( .OUT(na340_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na401_2), .IN7(1'b1), .IN8(na341_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x68y84     80'h00_0018_00_0000_0888_CCCD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a341_1 ( .OUT(na341_1), .IN1(~na374_1), .IN2(na343_1), .IN3(1'b0), .IN4(na378_1), .IN5(1'b0), .IN6(na396_1), .IN7(1'b0),
                     .IN8(na378_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x71y80     80'h00_0018_00_0000_0EEE_DDDE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(na358_1), .IN2(na346_1), .IN3(~na8371_1), .IN4(na406_1), .IN5(~na6816_2), .IN6(na346_2), .IN7(~na8371_2),
                     .IN8(na406_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x74y72     80'h00_0060_00_0000_0C08_FF23
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a344_4 ( .OUT(na344_2), .IN1(1'b1), .IN2(~na173_1), .IN3(na34_2), .IN4(~na5585_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x65y82     80'h00_0078_00_0000_0C88_4FA2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a346_1 ( .OUT(na346_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na347_1), .IN8(na48_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a346_4 ( .OUT(na346_2), .IN1(na5261_1), .IN2(~na9890_2), .IN3(na517_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y81     80'h00_0078_00_0000_0C88_114F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_1 ( .OUT(na347_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na348_1), .IN6(~na351_1), .IN7(~na350_1), .IN8(~na349_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a347_4 ( .OUT(na347_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na9217_2), .IN4(na48_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y83     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_1 ( .OUT(na348_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na50_2), .IN6(na3984_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y82     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3491_1), .IN8(na5695_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y83     80'h00_0018_00_0040_0A32_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a350_1 ( .OUT(na350_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3986_1), .IN6(~na3489_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y82     80'h00_0018_00_0040_0A51_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1377_1), .IN5(~na3487_1), .IN6(1'b0), .IN7(na5697_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////D      x65y73     80'h00_F618_00_0040_0C89_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1), .IN1(na356_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na6803_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1), .IN8(~na9911_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a353_5 ( .OUT(na353_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na353_1) );
// C_MX2b////D      x70y71     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6354_1), .IN8(na355_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a354_5 ( .OUT(na354_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na354_1) );
// C_MX4a////      x62y66     80'h00_0018_00_0040_0C06_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1), .IN1(1'b0), .IN2(na5957_2), .IN3(na5264_2), .IN4(1'b0), .IN5(na3264_1), .IN6(1'b1), .IN7(~na3265_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x65y65     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na357_1), .IN8(na6343_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a356_5 ( .OUT(na356_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na356_1) );
// C_MX4a////      x62y67     80'h00_0018_00_0040_0C06_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b0), .IN2(na5956_1), .IN3(na5263_1), .IN4(1'b0), .IN5(na3264_1), .IN6(1'b1), .IN7(~na3265_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x65y75     80'h00_0018_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1372_1), .IN6(na9247_2), .IN7(na359_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x66y81     80'h00_0078_00_0000_0C88_AA33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3262_1), .IN6(1'b1), .IN7(na517_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a359_4 ( .OUT(na359_2), .IN1(1'b1), .IN2(~na399_1), .IN3(1'b1), .IN4(~na404_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x69y73     80'h00_0060_00_0000_0C08_FFD3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a364_4 ( .OUT(na364_2), .IN1(1'b0), .IN2(~na2554_1), .IN3(~na2558_1), .IN4(na6810_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y70     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a365_4 ( .OUT(na365_2), .IN1(~na2565_1), .IN2(~na2564_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x61y72     80'h00_FA18_00_0000_0788_F3FC
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a369_1 ( .OUT(na369_1), .IN1(1'b1), .IN2(na2557_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2554_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a369_5 ( .OUT(na369_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na369_1) );
// C_ORAND////      x71y83     80'h00_0018_00_0000_0888_FCCE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_1 ( .OUT(na374_1), .IN1(na402_1), .IN2(na401_2), .IN3(1'b0), .IN4(na378_2), .IN5(1'b0), .IN6(na1462_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x72y92     80'h00_0078_00_0000_0C88_5331
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3610_2), .IN7(~na47_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a378_4 ( .OUT(na378_2), .IN1(~na1392_1), .IN2(~na9514_2), .IN3(1'b1), .IN4(~na1481_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x73y75     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_1 ( .OUT(na379_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2565_1), .IN6(~na2557_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x70y73     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a380_4 ( .OUT(na380_2), .IN1(~na2566_1), .IN2(na365_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y74     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a383_4 ( .OUT(na383_2), .IN1(na9617_2), .IN2(na2557_1), .IN3(na380_2), .IN4(na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x66y74     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a385_1 ( .OUT(na385_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2576_2), .IN6(~na2578_2), .IN7(~na9630_2),
                     .IN8(~na2582_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x76y75     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2562_1), .IN6(~na2561_1), .IN7(~na2560_1),
                     .IN8(~na2563_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y78     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a387_4 ( .OUT(na387_2), .IN1(~na2584_2), .IN2(~na2586_2), .IN3(na3307_2), .IN4(na389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x66y80     80'h00_0078_00_0000_0C88_1F22
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a389_1 ( .OUT(na389_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2588_2), .IN8(~na2590_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a389_4 ( .OUT(na389_2), .IN1(na2584_2), .IN2(~na2586_2), .IN3(na2588_2), .IN4(~na2590_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x70y74     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a393_4 ( .OUT(na393_2), .IN1(1'b1), .IN2(na2553_1), .IN3(na2552_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x67y84     80'h00_0018_00_0000_0888_7F3C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_1 ( .OUT(na396_1), .IN1(1'b0), .IN2(na397_2), .IN3(1'b0), .IN4(~na42_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na517_2), .IN8(~na3562_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y80     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a397_4 ( .OUT(na397_2), .IN1(1'b1), .IN2(na9205_2), .IN3(na8371_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y86     80'h00_0018_00_0000_0888_143C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b1), .IN2(na521_1), .IN3(1'b1), .IN4(~na404_2), .IN5(~na9511_2), .IN6(na505_2), .IN7(~na507_1),
                     .IN8(~na404_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x71y74     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a401_4 ( .OUT(na401_2_i), .IN1(na6823_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a401_5 ( .OUT(na401_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na401_2_i) );
// C_AND////      x73y85     80'h00_0018_00_0000_0C88_32FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a402_1 ( .OUT(na402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na712_1), .IN6(~na173_1), .IN7(1'b1), .IN8(~na9675_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////D      x72y89     80'h00_FE18_00_0000_0888_7F35
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1), .IN1(~na2994_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3200_1),
                     .IN8(~na2679_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a403_5 ( .OUT(na403_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na403_1) );
// C_AND/D//AND/D      x64y80     80'h00_FE00_80_0000_0C88_8F2A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a404_1 ( .OUT(na404_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na404_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a404_2 ( .OUT(na404_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na404_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a404_4 ( .OUT(na404_2_i), .IN1(na407_2), .IN2(1'b1), .IN3(na403_1), .IN4(~na406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a404_5 ( .OUT(na404_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na404_2_i) );
// C_AND///AND/      x64y74     80'h00_0078_00_0000_0C88_2484
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a406_1 ( .OUT(na406_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na5930_1), .IN6(na5977_1), .IN7(na517_2), .IN8(~na344_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a406_4 ( .OUT(na406_2), .IN1(~na353_1), .IN2(na3325_1), .IN3(na517_1), .IN4(na523_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x69y87     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a407_4 ( .OUT(na407_2), .IN1(1'b0), .IN2(na397_2), .IN3(na507_1), .IN4(na42_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x65y76     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1038_1), .IN6(1'b1), .IN7(na409_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a408_2 ( .OUT(na408_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na408_1_i) );
// C_AND////      x72y85     80'h00_0018_00_0000_0888_34CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a409_1 ( .OUT(na409_1), .IN1(na1126_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1864_2), .IN5(~na1126_1), .IN6(na410_1), .IN7(1'b1),
                     .IN8(~na1864_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x71y90     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a410_1 ( .OUT(na410_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(na1358_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x67y61     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a412_4 ( .OUT(na412_2_i), .IN1(na1038_2), .IN2(1'b1), .IN3(na409_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a412_5 ( .OUT(na412_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na412_2_i) );
// C_AND/D///      x53y74     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na878_1), .IN6(1'b1), .IN7(na409_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a413_2 ( .OUT(na413_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na413_1_i) );
// C_///AND/D      x59y68     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a414_4 ( .OUT(na414_2_i), .IN1(na878_2), .IN2(1'b1), .IN3(na409_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a414_5 ( .OUT(na414_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na414_2_i) );
// C_AND/D///      x56y85     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na409_1), .IN8(na984_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a415_2 ( .OUT(na415_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na415_1_i) );
// C_AND/D///      x78y60     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na409_1), .IN8(na984_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a416_2 ( .OUT(na416_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na416_1_i) );
// C_AND*/D///      x65y80     80'h00_F600_00_0000_0388_C3FF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a417_1 ( .OUT(na417_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na46_1), .IN7(1'b1), .IN8(na404_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a417_2 ( .OUT(na417_1), .CLK(na4116_1), .EN(~na359_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na417_1_i) );
// C_AND/D///      x58y83     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a418_1 ( .OUT(na418_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na409_1), .IN8(na999_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a418_2 ( .OUT(na418_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na418_1_i) );
// C_AND/D///      x57y75     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a419_1 ( .OUT(na419_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na409_1), .IN8(na999_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a419_2 ( .OUT(na419_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na419_1_i) );
// C_MX4b/D///      x90y71     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a420_1 ( .OUT(na420_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na420_1),
                     .IN8(na61_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a420_2 ( .OUT(na420_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na420_1_i) );
// C_ORAND////      x91y73     80'h00_0018_00_0000_0888_FDD5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(~na9184_2), .IN2(1'b0), .IN3(~na9187_2), .IN4(na154_1), .IN5(~na214_2), .IN6(na9179_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x89y65     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na66_1), .IN8(na9221_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_2 ( .OUT(na423_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na423_1_i) );
// C_MX4b/D///      x92y74     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a424_1 ( .OUT(na424_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na63_1), .IN8(na424_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a424_2 ( .OUT(na424_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na424_1_i) );
// C_MX4b/D///      x99y73     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1_i), .IN1(na426_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na425_1), .IN6(na259_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_2 ( .OUT(na425_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na425_1_i) );
// C_///AND/      x101y73     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a426_4 ( .OUT(na426_2), .IN1(na9229_2), .IN2(1'b1), .IN3(na427_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y75     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a427_4 ( .OUT(na427_2), .IN1(na9954_2), .IN2(~na435_1), .IN3(na433_1), .IN4(na9223_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y77     80'h00_0078_00_0000_0C88_8FA2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a428_1 ( .OUT(na428_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na430_1), .IN8(na429_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a428_4 ( .OUT(na428_2), .IN1(na9166_2), .IN2(~na89_1), .IN3(na8_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x102y82     80'h00_0060_00_0000_0C0E_FF5A
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a429_4 ( .OUT(na429_2), .IN1(na6828_1), .IN2(1'b0), .IN3(~na8_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x100y77     80'h00_0018_00_0000_0888_DF33
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_1 ( .OUT(na430_1), .IN1(1'b0), .IN2(~na431_1), .IN3(1'b0), .IN4(~na41_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na8_1), .IN8(na9225_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y76     80'h00_0018_00_0000_0888_FCEA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1), .IN1(na9_1), .IN2(1'b0), .IN3(na63_1), .IN4(na37_1), .IN5(1'b0), .IN6(na31_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y67     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a432_1 ( .OUT(na432_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na85_1), .IN7(~na84_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x94y77     80'h00_0078_00_0000_0C88_2A85
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a433_1 ( .OUT(na433_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na88_1), .IN6(1'b1), .IN7(na8_1), .IN8(~na87_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a433_4 ( .OUT(na433_2), .IN1(~na88_1), .IN2(1'b1), .IN3(na8_1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y82     80'h00_0078_00_0000_0C88_AC8A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na91_1), .IN7(na8_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a435_4 ( .OUT(na435_2), .IN1(na88_1), .IN2(1'b1), .IN3(na8_1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y79     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a436_1 ( .OUT(na436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na155_1), .IN6(1'b1), .IN7(na8_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x94y73     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na437_1),
                     .IN8(na37_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_2 ( .OUT(na437_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na437_1_i) );
// C_MX4b/D///      x93y65     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na438_1), .IN6(na35_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_2 ( .OUT(na438_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na438_1_i) );
// C_MX4b/D///      x88y63     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_1 ( .OUT(na439_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na439_1),
                     .IN8(na39_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_2 ( .OUT(na439_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na439_1_i) );
// C_MX4b/D///      x94y74     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_1 ( .OUT(na440_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na84_1), .IN8(na440_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_2 ( .OUT(na440_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na440_1_i) );
// C_MX4b/D///      x87y65     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a441_1 ( .OUT(na441_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na441_1), .IN6(na85_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a441_2 ( .OUT(na441_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na441_1_i) );
// C_MX4b/D///      x91y74     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na86_1), .IN6(na442_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_2 ( .OUT(na442_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na442_1_i) );
// C_MX4b/D///      x109y77     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1_i), .IN1(na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na443_1), .IN6(na6481_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_2 ( .OUT(na443_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na443_1_i) );
// C_AND////      x107y79     80'h00_0018_00_0000_0C88_C4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a444_1 ( .OUT(na444_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10027_2), .IN6(na2931_1), .IN7(1'b1), .IN8(na154_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x98y71     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a445_1 ( .OUT(na445_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na445_1),
                     .IN8(na87_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a445_2 ( .OUT(na445_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na445_1_i) );
// C_MX4b/D///      x93y70     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a446_1 ( .OUT(na446_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na88_1), .IN6(na446_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a446_2 ( .OUT(na446_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na446_1_i) );
// C_MX4b/D///      x103y85     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a447_1 ( .OUT(na447_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na447_1), .IN6(na454_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a447_2 ( .OUT(na447_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na447_1_i) );
// C_AND////      x105y81     80'h00_0018_00_0000_0888_2F23
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a448_1 ( .OUT(na448_1), .IN1(1'b1), .IN2(~na435_1), .IN3(na436_1), .IN4(~na452_1), .IN5(1'b1), .IN6(1'b1), .IN7(na8_2), .IN8(~na452_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y76     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2), .IN1(~na86_1), .IN2(~na9154_2), .IN3(na8_1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x98y86     80'h00_0078_00_0000_0C88_AEAE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na88_1), .IN6(na9161_2), .IN7(na8_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a452_4 ( .OUT(na452_2), .IN1(na9164_2), .IN2(na89_1), .IN3(na8_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x101y86     80'h00_0078_00_0000_0C88_5CAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a454_1 ( .OUT(na454_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a454_4 ( .OUT(na454_2), .IN1(na488_1), .IN2(1'b1), .IN3(na490_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x100y70     80'h00_FE00_00_0040_0AC3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1_i), .IN1(~na426_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na260_1),
                     .IN8(na455_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a455_2 ( .OUT(na455_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na455_1_i) );
// C_MX4b/D///      x89y73     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a456_1 ( .OUT(na456_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na90_1), .IN8(na9233_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a456_2 ( .OUT(na456_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na456_1_i) );
// C_MX4b/D///      x107y83     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_1 ( .OUT(na457_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9236_2),
                     .IN8(na9234_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_2 ( .OUT(na457_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na457_1_i) );
// C_AND////      x99y78     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a459_1 ( .OUT(na459_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(na435_2), .IN7(na436_1), .IN8(na9228_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y83     80'h00_0078_00_0000_0C88_4FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a463_1 ( .OUT(na463_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(na2536_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a463_4 ( .OUT(na463_2), .IN1(na428_1), .IN2(na459_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x93y69     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a464_1 ( .OUT(na464_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na464_1), .IN6(na91_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a464_2 ( .OUT(na464_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na464_1_i) );
// C_AND////      x83y74     80'h00_0018_00_0000_0888_8884
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1), .IN1(~na9140_2), .IN2(na12_1), .IN3(na469_1), .IN4(na28_1), .IN5(na19_1), .IN6(na13_1), .IN7(na469_2),
                     .IN8(na20_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y73     80'h00_0018_00_0000_0888_CC88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a468_1 ( .OUT(na468_1), .IN1(na19_1), .IN2(na13_1), .IN3(na469_2), .IN4(na20_1), .IN5(1'b1), .IN6(na12_1), .IN7(1'b1), .IN8(na28_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x82y73     80'h00_0078_00_0000_0C88_8A88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a469_1 ( .OUT(na469_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na29_1), .IN6(1'b1), .IN7(na30_1), .IN8(na21_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a469_4 ( .OUT(na469_2), .IN1(na17_1), .IN2(na15_1), .IN3(na9136_2), .IN4(na16_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x99y72     80'h00_FE00_00_0040_0A31_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na19_1), .IN6(na470_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_2 ( .OUT(na470_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na470_1_i) );
// C_MX4b/D///      x109y85     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_1 ( .OUT(na471_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na471_1), .IN6(na472_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_2 ( .OUT(na471_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na471_1_i) );
// C_AND////      x99y84     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a472_1 ( .OUT(na472_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na9404_2), .IN7(na2538_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x96y75     80'h00_FE00_00_0040_0AC8_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a473_1 ( .OUT(na473_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na473_1),
                     .IN8(~na20_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a473_2 ( .OUT(na473_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na473_1_i) );
// C_MX4b/D///      x101y77     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a474_1 ( .OUT(na474_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na474_1), .IN6(~na12_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a474_2 ( .OUT(na474_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na474_1_i) );
// C_MX4b/D///      x99y71     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_1 ( .OUT(na475_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na475_1), .IN6(~na13_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_2 ( .OUT(na475_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na475_1_i) );
// C_MX4b/D///      x91y71     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_1 ( .OUT(na476_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na476_1), .IN6(~na15_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_2 ( .OUT(na476_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na476_1_i) );
// C_MX4b/D///      x96y77     80'h00_FE00_00_0040_0AC8_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na477_1),
                     .IN8(~na16_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_2 ( .OUT(na477_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na477_1_i) );
// C_AND///AND/      x100y67     80'h00_0078_00_0000_0C88_C58F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a478_1 ( .OUT(na478_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9947_2), .IN6(1'b1), .IN7(1'b1), .IN8(na6673_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a478_4 ( .OUT(na478_2), .IN1(1'b1), .IN2(1'b1), .IN3(na8_1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y81     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a479_1 ( .OUT(na479_1_i), .IN1(1'b1), .IN2(na981_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na479_1), .IN6(na9863_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a479_2 ( .OUT(na479_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na479_1_i) );
// C_MX4b/D///      x109y79     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a480_1 ( .OUT(na480_1_i), .IN1(1'b1), .IN2(na981_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na480_1), .IN6(na4177_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a480_2 ( .OUT(na480_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na480_1_i) );
// C_MX4b/D///      x105y85     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a481_1 ( .OUT(na481_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na481_1), .IN6(na482_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a481_2 ( .OUT(na481_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na481_1_i) );
// C_///AND/      x97y86     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a482_4 ( .OUT(na482_2), .IN1(1'b1), .IN2(~na9404_2), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x105y86     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a483_1 ( .OUT(na483_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9236_2),
                     .IN8(na9238_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a483_2 ( .OUT(na483_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na483_1_i) );
// C_MX4b/D///      x95y79     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_1 ( .OUT(na484_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na484_1), .IN6(~na24_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_2 ( .OUT(na484_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na484_1_i) );
// C_MX4b/D///      x94y80     80'h00_FE00_00_0040_0AC4_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a485_1 ( .OUT(na485_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na22_1),
                     .IN8(na485_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a485_2 ( .OUT(na485_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na485_1_i) );
// C_MX4b/D///      x103y86     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9239_2), .IN6(na454_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_2 ( .OUT(na486_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na486_1_i) );
// C_AND///AND/      x105y77     80'h00_0078_00_0000_0C88_8231
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a488_1 ( .OUT(na488_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9947_2), .IN6(~na36_1), .IN7(na489_1), .IN8(na429_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a488_4 ( .OUT(na488_2), .IN1(~na854_1), .IN2(~na450_2), .IN3(1'b1), .IN4(~na429_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y79     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_1 ( .OUT(na489_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na432_1), .IN8(~na41_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y87     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a490_4 ( .OUT(na490_2), .IN1(na9954_2), .IN2(~na435_1), .IN3(na433_2), .IN4(na9230_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x94y79     80'h00_FE00_00_0040_0AC8_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a492_1 ( .OUT(na492_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na492_1),
                     .IN8(~na23_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a492_2 ( .OUT(na492_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na492_1_i) );
// C_MX4b/D///      x91y77     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_1 ( .OUT(na493_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na493_1), .IN6(~na25_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_2 ( .OUT(na493_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na493_1_i) );
// C_MX4b/D///      x93y79     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a494_1 ( .OUT(na494_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na494_1), .IN6(~na27_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a494_2 ( .OUT(na494_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na494_1_i) );
// C_MX4b/D///      x98y75     80'h00_FE00_00_0040_0AC8_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na495_1),
                     .IN8(~na28_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_2 ( .OUT(na495_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na495_1_i) );
// C_MX4b/D///      x93y78     80'h00_FE00_00_0040_0A31_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a496_1 ( .OUT(na496_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na29_1), .IN6(na496_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a496_2 ( .OUT(na496_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na496_1_i) );
// C_MX4b/D///      x98y80     80'h00_FE00_00_0040_0AC4_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_1 ( .OUT(na497_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na30_1),
                     .IN8(na497_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_2 ( .OUT(na497_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na497_1_i) );
// C_AND/D//AND/D      x130y47     80'h00_FE00_80_0000_0C88_CC4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a498_1 ( .OUT(na498_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3874_2), .IN7(1'b1), .IN8(na499_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a498_2 ( .OUT(na498_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na498_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a498_4 ( .OUT(na498_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na498_2), .IN4(na499_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a498_5 ( .OUT(na498_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na498_2_i) );
// C_///AND/      x126y56     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a499_4 ( .OUT(na499_2), .IN1(1'b1), .IN2(~na9941_2), .IN3(1'b1), .IN4(~na500_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x130y54     80'h00_FE18_00_0000_0888_558F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a500_1 ( .OUT(na500_1), .IN1(1'b1), .IN2(1'b1), .IN3(na498_1), .IN4(na3204_1), .IN5(~na790_2), .IN6(1'b1), .IN7(~na498_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a500_5 ( .OUT(na500_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na500_1) );
// C_ORAND/D///      x69y87     80'h00_FE00_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na501_1), .IN6(na504_1), .IN7(na502_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a501_2 ( .OUT(na501_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na501_1_i) );
// C_///AND/      x66y89     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a502_4 ( .OUT(na502_2), .IN1(na9214_2), .IN2(na521_1), .IN3(na1492_1), .IN4(na503_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x70y92     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a503_4 ( .OUT(na503_2), .IN1(1'b1), .IN2(na396_1), .IN3(1'b1), .IN4(na378_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x59y72     80'h00_0018_00_0000_0888_B335
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a504_1 ( .OUT(na504_1), .IN1(~na358_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na406_1), .IN5(1'b0), .IN6(~na9219_2), .IN7(na347_1),
                     .IN8(~na48_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x67y88     80'h00_FE00_80_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a505_1 ( .OUT(na505_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na502_2), .IN8(na6834_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a505_2 ( .OUT(na505_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na505_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a505_4 ( .OUT(na505_2_i), .IN1(1'b1), .IN2(na505_1), .IN3(na502_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a505_5 ( .OUT(na505_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na505_2_i) );
// C_///AND/      x69y84     80'h00_0060_00_0000_0C08_FF2C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a506_4 ( .OUT(na506_2), .IN1(1'b1), .IN2(na521_1), .IN3(na1492_1), .IN4(~na406_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x68y85     80'h00_FE00_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a507_1 ( .OUT(na507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6836_1), .IN6(na508_1), .IN7(na403_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a507_2 ( .OUT(na507_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na507_1_i) );
// C_AND////      x61y84     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a508_1 ( .OUT(na508_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na407_2), .IN6(1'b1), .IN7(1'b1), .IN8(na406_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x71y81     80'h00_0078_00_0000_0C88_3883
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a511_1 ( .OUT(na511_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9218_2), .IN6(na397_2), .IN7(1'b1), .IN8(~na42_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a511_4 ( .OUT(na511_2), .IN1(1'b1), .IN2(~na343_1), .IN3(na1492_1), .IN4(na503_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y83     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a514_4 ( .OUT(na514_2), .IN1(1'b1), .IN2(na396_1), .IN3(~na47_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x104y84     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a515_1 ( .OUT(na515_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6841_1), .IN6(na516_1), .IN7(1'b0), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a515_2 ( .OUT(na515_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na515_1_i) );
// C_AND////      x103y84     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a516_1 ( .OUT(na516_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2925_1), .IN6(1'b1), .IN7(na298_1), .IN8(na154_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND/D      x68y79     80'h00_FE00_80_0000_0C88_AEAE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a517_1 ( .OUT(na517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na511_2), .IN6(na6839_2), .IN7(na403_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a517_2 ( .OUT(na517_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na517_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a517_4 ( .OUT(na517_2_i), .IN1(na511_1), .IN2(na6839_1), .IN3(na403_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a517_5 ( .OUT(na517_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na517_2_i) );
// C_AND////D      x72y88     80'h00_FA18_00_0000_0888_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a520_1 ( .OUT(na520_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3259_1), .IN7(1'b1), .IN8(na1399_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a520_5 ( .OUT(na520_2), .CLK(na4116_1), .EN(na522_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na520_1) );
// C_ORAND/D///      x69y88     80'h00_FE00_00_0000_0888_AAE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a521_1 ( .OUT(na521_1_i), .IN1(1'b0), .IN2(~na399_1), .IN3(na6845_2), .IN4(na520_1), .IN5(na1388_1), .IN6(1'b0), .IN7(na403_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a521_2 ( .OUT(na521_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na521_1_i) );
// C_///ORAND/      x71y77     80'h00_0060_00_0000_0C08_FFEA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a522_4 ( .OUT(na522_2), .IN1(na1388_1), .IN2(1'b0), .IN3(na6845_2), .IN4(na520_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x72y74     80'h00_FE00_00_0000_0888_FDAD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1_i), .IN1(~na6847_1), .IN2(na9249_2), .IN3(na403_1), .IN4(1'b0), .IN5(~na9143_2), .IN6(na173_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a523_2 ( .OUT(na523_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na523_1_i) );
// C_///AND/      x61y81     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a526_4 ( .OUT(na526_2), .IN1(na9204_2), .IN2(na504_1), .IN3(na3308_1), .IN4(na3324_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x62y76     80'h00_0018_00_0040_0C4A_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a527_1 ( .OUT(na527_1), .IN1(1'b0), .IN2(na5953_1), .IN3(1'b1), .IN4(na9250_2), .IN5(1'b1), .IN6(na5953_2), .IN7(~na357_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x63y79     80'h00_0018_00_0000_0888_77D7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a528_1 ( .OUT(na528_1), .IN1(~na3313_1), .IN2(~na417_1), .IN3(~na531_2), .IN4(na6853_2), .IN5(~na3313_2), .IN6(~na9565_2),
                     .IN7(~na5456_1), .IN8(~na3309_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x72y87     80'h00_FE00_80_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a531_1 ( .OUT(na531_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na6855_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a531_2 ( .OUT(na531_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na531_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a531_4 ( .OUT(na531_2_i), .IN1(1'b1), .IN2(na6849_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a531_5 ( .OUT(na531_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na531_2_i) );
// C_MX4a////      x62y80     80'h00_0018_00_0040_0C4A_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a532_1 ( .OUT(na532_1), .IN1(1'b0), .IN2(na5953_1), .IN3(1'b1), .IN4(na9251_2), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1), .IN8(~na355_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x67y85     80'h00_0018_00_0000_0888_77D7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1), .IN1(~na3313_1), .IN2(~na640_2), .IN3(~na531_1), .IN4(na6859_1), .IN5(~na3313_2), .IN6(~na2173_1),
                     .IN7(~na5457_1), .IN8(~na3309_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////D      x55y78     80'h00_FA18_00_0040_0CB3_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a536_1 ( .OUT(na536_1), .IN1(~na537_1), .IN2(~na5953_1), .IN3(1'b0), .IN4(1'b1), .IN5(na540_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na9912_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a536_5 ( .OUT(na536_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na536_1) );
// C_ORAND////      x69y79     80'h00_0018_00_0000_0888_77B7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a537_1 ( .OUT(na537_1), .IN1(~na3313_1), .IN2(~na1125_2), .IN3(na6864_1), .IN4(~na9258_2), .IN5(~na3313_2), .IN6(~na2175_1),
                     .IN7(~na5458_2), .IN8(~na3309_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y71     80'h00_0018_00_0040_0A94_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a540_1 ( .OUT(na540_1), .IN1(1'b1), .IN2(~na9804_2), .IN3(~na9803_2), .IN4(1'b1), .IN5(na5958_1), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na5265_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////D      x68y87     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a542_1 ( .OUT(na542_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na3539_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na545_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a542_5 ( .OUT(na542_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na542_1) );
// C_MX4b////      x58y75     80'h00_0018_00_0040_0A60_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a545_1 ( .OUT(na545_1), .IN1(1'b1), .IN2(na9804_2), .IN3(~na9803_2), .IN4(1'b1), .IN5(1'b0), .IN6(na5959_2), .IN7(na9891_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x73y87     80'h00_FE00_80_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a546_1 ( .OUT(na546_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6871_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a546_2 ( .OUT(na546_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na546_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a546_4 ( .OUT(na546_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na6866_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a546_5 ( .OUT(na546_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na546_2_i) );
// C_MX4a////D      x68y74     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a547_1 ( .OUT(na547_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na548_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na550_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a547_5 ( .OUT(na547_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na547_1) );
// C_ORAND////      x58y82     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a548_1 ( .OUT(na548_1), .IN1(~na3313_2), .IN2(~na2179_1), .IN3(~na5460_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na551_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x62y69     80'h00_0018_00_0040_0A60_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a550_1 ( .OUT(na550_1), .IN1(1'b1), .IN2(na9804_2), .IN3(~na9803_2), .IN4(1'b1), .IN5(1'b0), .IN6(na5960_1), .IN7(na9892_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x66y84     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a551_1 ( .OUT(na551_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6875_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a551_2 ( .OUT(na551_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na551_1_i) );
// C_MX4a////D      x56y82     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a552_1 ( .OUT(na552_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na555_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na2369_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a552_5 ( .OUT(na552_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na552_1) );
// C_///AND/      x59y69     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a554_4 ( .OUT(na554_2), .IN1(~na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x62y84     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a555_1 ( .OUT(na555_1), .IN1(~na3313_2), .IN2(~na2181_1), .IN3(~na5461_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na557_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x70y90     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a557_4 ( .OUT(na557_2_i), .IN1(1'b1), .IN2(na6879_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a557_5 ( .OUT(na557_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na557_2_i) );
// C_MX4b/D///      x95y83     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a558_1 ( .OUT(na558_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na558_1), .IN6(na472_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a558_2 ( .OUT(na558_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na558_1_i) );
// C_MX4b/D///      x99y92     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a560_1 ( .OUT(na560_1_i), .IN1(~na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na5185_2), .IN6(na560_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a560_2 ( .OUT(na560_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na560_1_i) );
// C_ORAND/D//AND/D      x96y85     80'h00_FE00_80_0000_0C88_3E8F
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a561_1 ( .OUT(na561_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6881_2), .IN6(na562_2), .IN7(1'b0), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a561_2 ( .OUT(na561_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na561_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a561_4 ( .OUT(na561_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na561_1), .IN4(na1346_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a561_5 ( .OUT(na561_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na561_2_i) );
// C_///ORAND/      x97y88     80'h00_0060_00_0000_0C08_FFA7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a562_4 ( .OUT(na562_2), .IN1(~na563_1), .IN2(~na1351_1), .IN3(na561_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x97y81     80'h00_FE00_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a563_1 ( .OUT(na563_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na564_1), .IN7(na567_1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a563_2 ( .OUT(na563_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na563_1_i) );
// C_AND////      x101y88     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a564_1 ( .OUT(na564_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na565_2), .IN7(na436_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y76     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a565_4 ( .OUT(na565_2), .IN1(na566_1), .IN2(na435_1), .IN3(na433_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y75     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a566_1 ( .OUT(na566_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9166_2), .IN6(na89_1), .IN7(na8_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y85     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9947_2), .IN6(na450_2), .IN7(na489_1), .IN8(~na9146_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x100y85     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a568_1 ( .OUT(na568_1_i), .IN1(na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na568_1),
                     .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a568_2 ( .OUT(na568_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na568_1_i) );
// C_///AND/      x95y87     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a569_4 ( .OUT(na569_2), .IN1(na428_1), .IN2(na564_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y86     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a570_1 ( .OUT(na570_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3042_1),
                     .IN8(na9267_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a570_2 ( .OUT(na570_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na570_1_i) );
// C_MX4b/D///      x103y75     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a571_1 ( .OUT(na571_1_i), .IN1(na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na571_1), .IN6(na6483_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a571_2 ( .OUT(na571_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na571_1_i) );
// C_AND////      x109y75     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a572_1 ( .OUT(na572_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8107_2), .IN6(1'b1), .IN7(na2950_1), .IN8(na2948_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x101y78     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a573_1 ( .OUT(na573_1_i), .IN1(~na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6480_1), .IN6(na573_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a573_2 ( .OUT(na573_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na573_1_i) );
// C_MX4a////D      x56y72     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a574_1 ( .OUT(na574_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na576_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na2348_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a574_5 ( .OUT(na574_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na574_1) );
// C_ORAND////      x58y88     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a576_1 ( .OUT(na576_1), .IN1(~na3313_2), .IN2(~na2183_1), .IN3(~na5462_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na578_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x66y88     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a578_1 ( .OUT(na578_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6886_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a578_2 ( .OUT(na578_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na578_1_i) );
// C_MX4b/D///      x104y86     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_1 ( .OUT(na579_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na581_1), .IN6(na9270_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_2 ( .OUT(na579_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na579_1_i) );
// C_AND///AND/      x103y87     80'h00_0078_00_0000_0C88_5AAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_1 ( .OUT(na581_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2537_1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a581_4 ( .OUT(na581_2), .IN1(1'b1), .IN2(na459_1), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////D      x59y82     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a582_1 ( .OUT(na582_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na584_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na9568_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a582_5 ( .OUT(na582_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na582_1) );
// C_AND////      x58y84     80'h00_0018_00_0000_0888_345C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a584_1 ( .OUT(na584_1), .IN1(1'b1), .IN2(na6888_1), .IN3(~na6887_1), .IN4(1'b1), .IN5(~na6891_2), .IN6(na6888_2), .IN7(1'b1),
                     .IN8(~na6889_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x68y86     80'h00_FE00_80_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_1 ( .OUT(na587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na6892_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a587_2 ( .OUT(na587_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na587_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a587_4 ( .OUT(na587_2_i), .IN1(na9216_2), .IN2(1'b1), .IN3(na7207_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a587_5 ( .OUT(na587_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na587_2_i) );
// C_MX4a////D      x72y72     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a588_1 ( .OUT(na588_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na9276_2), .IN5(1'b1), .IN6(na5953_2), .IN7(~na589_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a588_5 ( .OUT(na588_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na588_1) );
// C_AND///AND/      x56y71     80'h00_0078_00_0000_0C88_CAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a589_1 ( .OUT(na589_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na554_2), .IN6(1'b1), .IN7(1'b1), .IN8(na5271_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a589_4 ( .OUT(na589_2), .IN1(1'b1), .IN2(na7905_2), .IN3(na2324_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y79     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a590_1 ( .OUT(na590_1), .IN1(~na3313_2), .IN2(~na2187_1), .IN3(~na5464_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na592_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x66y84     80'h00_FE00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a592_4 ( .OUT(na592_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na6896_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a592_5 ( .OUT(na592_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na592_2_i) );
// C_MX4a////D      x62y74     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a593_1 ( .OUT(na593_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na595_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na594_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a593_5 ( .OUT(na593_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na593_1) );
// C_AND////      x68y72     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_1 ( .OUT(na594_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na554_2), .IN6(na5272_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x64y78     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a595_1 ( .OUT(na595_1), .IN1(~na3313_2), .IN2(~na2189_1), .IN3(~na5465_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na597_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x66y82     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a597_1 ( .OUT(na597_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na6900_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a597_2 ( .OUT(na597_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na597_1_i) );
// C_MX4a////D      x62y70     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a598_1 ( .OUT(na598_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na600_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na2327_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a598_5 ( .OUT(na598_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na598_1) );
// C_ORAND////      x58y86     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a600_1 ( .OUT(na600_1), .IN1(~na3313_2), .IN2(~na2191_1), .IN3(~na5466_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na602_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x68y80     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a602_4 ( .OUT(na602_2_i), .IN1(na9216_2), .IN2(1'b1), .IN3(na6904_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a602_5 ( .OUT(na602_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na602_2_i) );
// C_MX4a////D      x60y74     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a603_1 ( .OUT(na603_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na604_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na607_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a603_5 ( .OUT(na603_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na603_1) );
// C_ORAND////      x70y82     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a604_1 ( .OUT(na604_1), .IN1(~na3313_2), .IN2(~na2195_1), .IN3(~na5468_1), .IN4(~na3309_1), .IN5(~na1405_1), .IN6(~na9816_2),
                     .IN7(~na3308_1), .IN8(~na9282_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y73     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a607_1 ( .OUT(na607_1), .IN1(na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na9893_2), .IN6(na5953_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x66y89     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a608_1 ( .OUT(na608_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6909_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a608_2 ( .OUT(na608_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na608_1_i) );
// C_MX4a////D      x58y80     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a609_1 ( .OUT(na609_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na610_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na612_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a609_5 ( .OUT(na609_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na609_1) );
// C_ORAND////      x62y82     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a610_1 ( .OUT(na610_1), .IN1(~na3313_2), .IN2(~na2197_1), .IN3(~na5469_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na613_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y72     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a612_1 ( .OUT(na612_1), .IN1(na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na9894_2), .IN6(na5953_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x66y88     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a613_4 ( .OUT(na613_2_i), .IN1(na6913_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a613_5 ( .OUT(na613_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na613_2_i) );
// C_MX4a////D      x56y84     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a614_1 ( .OUT(na614_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na615_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na617_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a614_5 ( .OUT(na614_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na614_1) );
// C_ORAND////      x62y90     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a615_1 ( .OUT(na615_1), .IN1(~na3313_2), .IN2(~na2201_1), .IN3(~na5471_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na618_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x58y76     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a617_1 ( .OUT(na617_1), .IN1(na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na9896_2), .IN6(na5956_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x70y84     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a618_1 ( .OUT(na618_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6917_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a618_2 ( .OUT(na618_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na618_1_i) );
// C_MX4a////D      x56y108     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a619_1 ( .OUT(na619_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na9289_2), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na622_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a619_5 ( .OUT(na619_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na619_1) );
// C_ORAND////      x57y89     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a620_1 ( .OUT(na620_1), .IN1(~na3313_2), .IN2(~na2199_1), .IN3(~na5470_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na623_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y76     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a622_1 ( .OUT(na622_1), .IN1(na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9895_2),
                     .IN8(na5955_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x70y88     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a623_4 ( .OUT(na623_2_i), .IN1(na6921_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a623_5 ( .OUT(na623_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na623_2_i) );
// C_MX4a////D      x54y102     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a624_1 ( .OUT(na624_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na625_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na627_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a624_5 ( .OUT(na624_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na624_1) );
// C_ORAND////      x62y86     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a625_1 ( .OUT(na625_1), .IN1(~na3313_2), .IN2(~na2203_1), .IN3(~na5472_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na628_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x58y77     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a627_1 ( .OUT(na627_1), .IN1(na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na9897_2), .IN6(na5957_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x70y92     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a628_1 ( .OUT(na628_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6925_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a628_2 ( .OUT(na628_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na628_1_i) );
// C_MX4a////D      x56y102     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a629_1 ( .OUT(na629_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na630_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na632_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a629_5 ( .OUT(na629_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na629_1) );
// C_ORAND////      x68y110     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a630_1 ( .OUT(na630_1), .IN1(~na3313_2), .IN2(~na2207_1), .IN3(~na5474_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na633_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x54y77     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a632_1 ( .OUT(na632_1), .IN1(na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na9898_2), .IN6(na5959_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x70y84     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a633_4 ( .OUT(na633_2_i), .IN1(na6929_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a633_5 ( .OUT(na633_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na633_2_i) );
// C_MX4a////D      x52y104     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a634_1 ( .OUT(na634_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na635_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na637_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a634_5 ( .OUT(na634_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na634_1) );
// C_ORAND////      x58y114     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1), .IN1(~na3313_2), .IN2(~na2209_1), .IN3(~na5475_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na638_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y73     80'h00_0018_00_0040_0AA0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a637_1 ( .OUT(na637_1), .IN1(1'b1), .IN2(~na9804_2), .IN3(~na9803_2), .IN4(1'b1), .IN5(1'b0), .IN6(na5960_1), .IN7(1'b0),
                     .IN8(na9899_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x70y90     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a638_1 ( .OUT(na638_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6933_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a638_2 ( .OUT(na638_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na638_1_i) );
// C_MX4b/D///      x105y88     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_1 ( .OUT(na639_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3044_1), .IN6(na639_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_2 ( .OUT(na639_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na639_1_i) );
// C_///AND*/D      x71y84     80'h00_F600_80_0000_0C07_FFC3
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a640_4 ( .OUT(na640_2_i), .IN1(1'b1), .IN2(~na1626_2), .IN3(1'b1), .IN4(na404_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a640_5 ( .OUT(na640_2), .CLK(na4116_1), .EN(~na359_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na640_2_i) );
// C_MX4b/D///      x107y82     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_1 ( .OUT(na641_1_i), .IN1(~na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6480_1), .IN6(na641_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_2 ( .OUT(na641_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na641_1_i) );
// C_AND////      x121y93     80'h00_0018_00_0000_0888_C1F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a643_1 ( .OUT(na643_1), .IN1(~na6936_2), .IN2(~na6937_2), .IN3(1'b1), .IN4(1'b1), .IN5(~na6936_1), .IN6(~na215_1), .IN7(1'b1),
                     .IN8(na654_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y98     80'h00_0018_00_0000_0888_8281
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a647_1 ( .OUT(na647_1), .IN1(~na7054_2), .IN2(~na6778_1), .IN3(na220_1), .IN4(na753_2), .IN5(na6776_1), .IN6(~na6778_2),
                     .IN7(na6777_2), .IN8(na6779_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y88     80'h00_0060_00_0000_0C08_FF84
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a649_4 ( .OUT(na649_2), .IN1(~na650_1), .IN2(na2894_2), .IN3(na2838_1), .IN4(na2836_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y87     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a650_1 ( .OUT(na650_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na652_2), .IN6(na9297_2), .IN7(na709_2), .IN8(~na753_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x125y97     80'h00_0078_00_0000_0C88_1F11
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a652_1 ( .OUT(na652_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na755_2), .IN8(~na753_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a652_4 ( .OUT(na652_2), .IN1(~na2951_2), .IN2(~na9719_2), .IN3(~na709_1), .IN4(~na2953_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x124y96     80'h00_0018_00_0000_0CEE_5A00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a654_1 ( .OUT(na654_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na6938_1), .IN6(1'b0), .IN7(~na2838_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y80     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2920_2), .IN6(1'b1), .IN7(1'b1), .IN8(na174_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x114y77     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a656_1 ( .OUT(na656_1), .IN1(1'b1), .IN2(na9169_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na102_1), .IN8(na92_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x125y98     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a657_1 ( .OUT(na657_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3737_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na654_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////D      x58y102     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a658_1 ( .OUT(na658_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na659_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na661_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a658_5 ( .OUT(na658_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na658_1) );
// C_ORAND////      x66y112     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a659_1 ( .OUT(na659_1), .IN1(~na3313_2), .IN2(~na2213_1), .IN3(~na5477_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na662_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y67     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a661_1 ( .OUT(na661_1), .IN1(na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9901_2),
                     .IN8(na5962_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x68y94     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a662_4 ( .OUT(na662_2_i), .IN1(1'b1), .IN2(na6942_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a662_5 ( .OUT(na662_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na662_2_i) );
// C_MX4b/D///      x110y86     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a663_1 ( .OUT(na663_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9236_2),
                     .IN8(na663_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a663_2 ( .OUT(na663_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na663_1_i) );
// C_MX4a////D      x62y108     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a664_1 ( .OUT(na664_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na665_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na667_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a664_5 ( .OUT(na664_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na664_1) );
// C_ORAND////      x66y116     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a665_1 ( .OUT(na665_1), .IN1(~na3313_2), .IN2(~na2215_1), .IN3(~na5478_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na668_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x58y74     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a667_1 ( .OUT(na667_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na5963_1), .IN6(na5285_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x74y86     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a668_1 ( .OUT(na668_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6946_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a668_2 ( .OUT(na668_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na668_1_i) );
// C_MX4a////D      x60y78     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a669_1 ( .OUT(na669_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na670_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na672_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a669_5 ( .OUT(na669_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na669_1) );
// C_ORAND////      x62y112     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a670_1 ( .OUT(na670_1), .IN1(~na3313_2), .IN2(~na2217_1), .IN3(~na5479_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na673_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x60y73     80'h00_0018_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a672_1 ( .OUT(na672_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na5964_1),
                     .IN8(na5286_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x68y88     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a673_4 ( .OUT(na673_2_i), .IN1(na6950_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a673_5 ( .OUT(na673_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na673_2_i) );
// C_MX4a////D      x58y106     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a674_1 ( .OUT(na674_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na675_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na677_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a674_5 ( .OUT(na674_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na674_1) );
// C_ORAND////      x62y114     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a675_1 ( .OUT(na675_1), .IN1(~na3313_2), .IN2(~na2219_1), .IN3(~na5480_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na678_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x60y77     80'h00_0018_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a677_1 ( .OUT(na677_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na5965_1),
                     .IN8(na5287_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x70y88     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a678_1 ( .OUT(na678_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6954_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a678_2 ( .OUT(na678_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na678_1_i) );
// C_MX4a////D      x56y104     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a679_1 ( .OUT(na679_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na680_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na682_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a679_5 ( .OUT(na679_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na679_1) );
// C_ORAND////      x64y114     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a680_1 ( .OUT(na680_1), .IN1(~na3313_2), .IN2(~na2221_1), .IN3(~na5481_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na683_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y74     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a682_1 ( .OUT(na682_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na5967_2), .IN6(na5288_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x70y86     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a683_4 ( .OUT(na683_2_i), .IN1(1'b1), .IN2(na6958_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a683_5 ( .OUT(na683_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na683_2_i) );
// C_MX4a////D      x60y108     80'h00_FA18_00_0040_0CB3_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a684_1 ( .OUT(na684_1), .IN1(~na685_1), .IN2(~na5953_1), .IN3(1'b0), .IN4(1'b1), .IN5(na687_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na9912_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a684_5 ( .OUT(na684_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na684_1) );
// C_ORAND////      x65y117     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1), .IN1(~na3313_2), .IN2(~na2223_1), .IN3(~na5482_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na688_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x67y67     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a687_1 ( .OUT(na687_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na5967_1), .IN6(na5289_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x66y92     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a688_1 ( .OUT(na688_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na6962_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a688_2 ( .OUT(na688_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na688_1_i) );
// C_MX4a////D      x56y106     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a689_1 ( .OUT(na689_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na690_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na692_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a689_5 ( .OUT(na689_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na689_1) );
// C_ORAND////      x60y118     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a690_1 ( .OUT(na690_1), .IN1(~na3313_2), .IN2(~na2225_1), .IN3(~na5483_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na693_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y75     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a692_1 ( .OUT(na692_1), .IN1(na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9902_2),
                     .IN8(na5969_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x66y82     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a693_4 ( .OUT(na693_2_i), .IN1(na6966_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a693_5 ( .OUT(na693_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na693_2_i) );
// C_MX4a////D      x62y102     80'h00_FA18_00_0040_0CB3_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a694_1 ( .OUT(na694_1), .IN1(~na695_1), .IN2(~na5953_1), .IN3(1'b0), .IN4(1'b1), .IN5(na697_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na9912_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a694_5 ( .OUT(na694_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na694_1) );
// C_ORAND////      x63y115     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1), .IN1(~na3313_2), .IN2(~na2227_1), .IN3(~na5484_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na698_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y67     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a697_1 ( .OUT(na697_1), .IN1(na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9903_2),
                     .IN8(na5969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x68y94     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a698_1 ( .OUT(na698_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6970_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a698_2 ( .OUT(na698_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na698_1_i) );
// C_MX4a////D      x64y108     80'h00_FA18_00_0040_0CBA_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a699_1 ( .OUT(na699_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na700_1), .IN5(1'b1), .IN6(na5953_2), .IN7(1'b1),
                     .IN8(~na702_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a699_5 ( .OUT(na699_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na699_1) );
// C_ORAND////      x66y114     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a700_1 ( .OUT(na700_1), .IN1(~na3313_2), .IN2(~na2229_1), .IN3(~na5485_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na703_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x62y78     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na5971_2), .IN6(na5292_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x68y90     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a703_4 ( .OUT(na703_2_i), .IN1(1'b1), .IN2(na6974_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a703_5 ( .OUT(na703_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na703_2_i) );
// C_MX4a////D      x60y80     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a704_1 ( .OUT(na704_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na705_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na707_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a704_5 ( .OUT(na704_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na704_1) );
// C_ORAND////      x68y116     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a705_1 ( .OUT(na705_1), .IN1(~na3313_2), .IN2(~na2231_1), .IN3(~na5486_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                     .IN8(~na708_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x60y75     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na5971_1), .IN6(na5293_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x68y92     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a708_4 ( .OUT(na708_2_i), .IN1(1'b1), .IN2(na6978_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a708_5 ( .OUT(na708_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na708_2_i) );
// C_ORAND/D//ORAND/D      x122y95     80'h00_FE00_80_0000_0C88_3E3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na710_1), .IN6(na6980_1), .IN7(1'b0), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_2 ( .OUT(na709_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na709_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a709_4 ( .OUT(na709_2_i), .IN1(na736_2), .IN2(na6995_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a709_5 ( .OUT(na709_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na709_2_i) );
// C_AND////      x129y97     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a710_1 ( .OUT(na710_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3735_2), .IN7(1'b1), .IN8(~na654_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x71y85     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na712_1), .IN6(1'b1), .IN7(~na9213_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x77y87     80'h00_FE00_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a712_1 ( .OUT(na712_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na711_1), .IN6(na713_1), .IN7(na403_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a712_2 ( .OUT(na712_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na712_1_i) );
// C_AND////      x71y96     80'h00_0018_00_0000_0888_54A1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a713_1 ( .OUT(na713_1), .IN1(~na711_1), .IN2(~na716_1), .IN3(na718_2), .IN4(1'b1), .IN5(~na714_2), .IN6(na9320_2), .IN7(~na718_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x71y91     80'h00_0078_00_0000_0C88_B3EC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a714_1 ( .OUT(na714_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na343_1), .IN7(na9208_2), .IN8(~na9513_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a714_4 ( .OUT(na714_2), .IN1(1'b0), .IN2(na396_1), .IN3(na47_2), .IN4(na9512_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x71y84     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a716_1 ( .OUT(na716_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na514_2), .IN6(1'b0), .IN7(na1408_1), .IN8(na9833_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x70y97     80'h00_0078_00_0000_0C88_8C24
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a718_1 ( .OUT(na718_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1414_2), .IN7(na1433_2), .IN8(na9509_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a718_4 ( .OUT(na718_2), .IN1(~na407_2), .IN2(na397_2), .IN3(na403_2), .IN4(~na404_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////D      x62y100     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na720_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na723_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a719_5 ( .OUT(na719_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na719_1) );
// C_ORAND////      x60y114     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a720_1 ( .OUT(na720_1), .IN1(~na3313_1), .IN2(~na5518_2), .IN3(~na5487_1), .IN4(~na3309_1), .IN5(~na3313_2), .IN6(~na2233_1),
                     .IN7(~na3308_1), .IN8(~na724_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x62y77     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na5972_1), .IN6(na5294_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x68y92     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a724_1 ( .OUT(na724_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6988_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a724_2 ( .OUT(na724_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na724_1_i) );
// C_ORAND/D///      x78y98     80'h00_FE00_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a725_1 ( .OUT(na725_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6990_1), .IN6(na713_1), .IN7(na403_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a725_2 ( .OUT(na725_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na725_1_i) );
// C_///ORAND/      x73y90     80'h00_0060_00_0000_0C08_FF7C
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a727_4 ( .OUT(na727_2), .IN1(1'b0), .IN2(na397_2), .IN3(~na517_2), .IN4(~na3562_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x75y88     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a728_1 ( .OUT(na728_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3909_1), .IN8(~na729_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a728_5 ( .OUT(na728_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na728_1) );
// C_MX2b////      x76y96     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a729_1 ( .OUT(na729_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3961_1), .IN8(na730_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x60y106     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a730_1 ( .OUT(na730_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2175_1), .IN7(1'b0), .IN8(~na9252_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x58y90     80'h00_0018_00_0000_0888_2ACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1), .IN1(na1372_1), .IN2(1'b1), .IN3(1'b1), .IN4(na5435_2), .IN5(na5927_1), .IN6(1'b1), .IN7(na5926_2),
                     .IN8(~na5435_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x71y87     80'h00_0060_00_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a734_4 ( .OUT(na734_2), .IN1(na714_1), .IN2(~na727_2), .IN3(na403_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y95     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a736_4 ( .OUT(na736_2), .IN1(1'b1), .IN2(na3735_1), .IN3(1'b1), .IN4(~na654_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x77y84     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3909_2), .IN8(~na738_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a737_5 ( .OUT(na737_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na737_1) );
// C_MX2b////      x74y98     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a738_1 ( .OUT(na738_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na739_1), .IN8(~na3964_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y113     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na731_1), .IN5(~na2177_1), .IN6(1'b0), .IN7(~na542_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x69y93     80'h00_FE00_80_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a740_1 ( .OUT(na740_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6996_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a740_2 ( .OUT(na740_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na740_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a740_4 ( .OUT(na740_2_i), .IN1(na6992_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a740_5 ( .OUT(na740_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na740_2_i) );
// C_MX2b////D      x73y89     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a741_1 ( .OUT(na741_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na742_1), .IN8(na3931_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a741_5 ( .OUT(na741_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na741_1) );
// C_MX2b////      x74y91     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a742_1 ( .OUT(na742_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3965_1), .IN8(na743_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y106     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a743_1 ( .OUT(na743_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2179_1), .IN7(1'b0), .IN8(~na547_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x75y95     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a745_1 ( .OUT(na745_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na746_1), .IN8(na3931_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a745_5 ( .OUT(na745_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na745_1) );
// C_MX2b////      x70y93     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a746_1 ( .OUT(na746_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na747_1), .IN8(~na3966_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y103     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a747_1 ( .OUT(na747_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2181_1), .IN7(1'b0), .IN8(~na552_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x69y94     80'h00_FE00_80_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a748_1 ( .OUT(na748_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6998_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a748_2 ( .OUT(na748_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na748_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a748_4 ( .OUT(na748_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na6997_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a748_5 ( .OUT(na748_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na748_2_i) );
// C_MX2b////D      x75y83     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a749_1 ( .OUT(na749_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3933_1), .IN8(~na750_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a749_5 ( .OUT(na749_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na749_1) );
// C_MX2b////      x74y84     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a750_1 ( .OUT(na750_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na5830_2), .IN6(na751_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y108     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a751_1 ( .OUT(na751_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2183_1), .IN7(1'b0), .IN8(~na574_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND/D      x120y94     80'h00_FE00_80_0000_0C88_3E3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_1 ( .OUT(na753_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7001_1), .IN6(na754_1), .IN7(1'b0), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_2 ( .OUT(na753_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na753_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a753_4 ( .OUT(na753_2_i), .IN1(na8113_1), .IN2(na2959_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a753_5 ( .OUT(na753_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na753_2_i) );
// C_AND////      x127y98     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a754_1 ( .OUT(na754_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3733_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na654_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x124y95     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a755_4 ( .OUT(na755_2_i), .IN1(na756_1), .IN2(na7003_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a755_5 ( .OUT(na755_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na755_2_i) );
// C_AND////      x125y95     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a756_1 ( .OUT(na756_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3733_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na654_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x94y85     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a757_1 ( .OUT(na757_1_i), .IN1(1'b1), .IN2(na758_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na757_1),
                     .IN8(na9330_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a757_2 ( .OUT(na757_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na757_1_i) );
// C_AND///AND/      x99y88     80'h00_0078_00_0000_0C88_AAA5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a758_1 ( .OUT(na758_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7004_2), .IN6(1'b1), .IN7(na3871_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a758_4 ( .OUT(na758_2), .IN1(~na7054_2), .IN2(1'b1), .IN3(na102_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x65y96     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_1 ( .OUT(na759_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na760_1), .IN8(na3935_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a759_5 ( .OUT(na759_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na759_1) );
// C_MX2b////      x76y81     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a760_1 ( .OUT(na760_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na5832_1), .IN6(na761_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y108     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a761_1 ( .OUT(na761_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2187_1), .IN7(1'b0), .IN8(~na588_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x73y82     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a763_1 ( .OUT(na763_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na764_1), .IN8(na3935_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a763_5 ( .OUT(na763_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na763_1) );
// C_MX2b////      x66y97     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a764_1 ( .OUT(na764_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na765_1), .IN8(~na3970_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y101     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2189_1), .IN7(1'b0), .IN8(~na593_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x69y95     80'h00_FE00_80_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a766_1 ( .OUT(na766_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na7007_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a766_2 ( .OUT(na766_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na766_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a766_4 ( .OUT(na766_2_i), .IN1(1'b1), .IN2(na7006_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a766_5 ( .OUT(na766_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na766_2_i) );
// C_MX2b////D      x76y92     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a767_1 ( .OUT(na767_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3937_1), .IN8(~na768_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a767_5 ( .OUT(na767_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na767_1) );
// C_MX2b////      x72y80     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a768_1 ( .OUT(na768_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b0), .IN4(1'b0), .IN5(na769_1), .IN6(~na5834_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y109     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a769_1 ( .OUT(na769_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2191_1), .IN7(1'b0), .IN8(~na598_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x62y92     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a771_1 ( .OUT(na771_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3937_2), .IN8(~na772_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a771_5 ( .OUT(na771_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na771_1) );
// C_MX2b////      x68y104     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a772_1 ( .OUT(na772_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3941_1), .IN8(na773_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y110     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a773_1 ( .OUT(na773_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na731_1), .IN5(1'b0), .IN6(~na1393_2), .IN7(1'b0), .IN8(~na2193_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x72y93     80'h00_FE00_80_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a774_1 ( .OUT(na774_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7009_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a774_2 ( .OUT(na774_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na774_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a774_4 ( .OUT(na774_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na7008_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a774_5 ( .OUT(na774_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na774_2_i) );
// C_MX2b////D      x74y88     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na776_1), .IN8(na3910_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a775_5 ( .OUT(na775_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na775_1) );
// C_MX2b////      x70y109     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a776_1 ( .OUT(na776_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na5836_2), .IN8(na777_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y116     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2195_1), .IN7(1'b0), .IN8(~na603_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x74y90     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na780_1), .IN8(na3910_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a779_5 ( .OUT(na779_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na779_1) );
// C_MX2b////      x70y99     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a780_1 ( .OUT(na780_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na781_1), .IN8(~na3943_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y105     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2197_1), .IN7(1'b0), .IN8(~na609_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x68y93     80'h00_FE00_80_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a782_1 ( .OUT(na782_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7011_1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a782_2 ( .OUT(na782_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na782_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a782_4 ( .OUT(na782_2_i), .IN1(na7010_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a782_5 ( .OUT(na782_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na782_2_i) );
// C_MX4b/D///      x94y84     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1_i), .IN1(1'b1), .IN2(~na758_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na784_2),
                     .IN8(na783_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_2 ( .OUT(na783_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na783_1_i) );
// C_///AND/      x98y83     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a784_4 ( .OUT(na784_2), .IN1(na7004_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na783_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x107y88     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_1 ( .OUT(na785_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9334_2), .IN6(na3046_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_2 ( .OUT(na785_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na785_1_i) );
// C_MX2b////D      x77y92     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a786_1 ( .OUT(na786_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3912_1), .IN8(~na787_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a786_5 ( .OUT(na786_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na786_1) );
// C_MX2b////      x76y84     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na5838_1), .IN8(na788_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x60y116     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a788_1 ( .OUT(na788_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2199_1), .IN7(1'b0), .IN8(~na619_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x131y47     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a790_4 ( .OUT(na790_2_i), .IN1(1'b1), .IN2(na3874_1), .IN3(1'b1), .IN4(na499_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a790_5 ( .OUT(na790_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na790_2_i) );
// C_MX4b/D///      x110y85     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_1 ( .OUT(na791_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9335_2), .IN6(na482_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_2 ( .OUT(na791_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na791_1_i) );
// C_MX2b////D      x75y90     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a792_1 ( .OUT(na792_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3912_2), .IN8(~na793_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a792_5 ( .OUT(na792_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na792_1) );
// C_MX2b////      x66y98     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a793_1 ( .OUT(na793_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3945_1), .IN8(na794_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y106     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a794_1 ( .OUT(na794_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2201_1), .IN7(1'b0), .IN8(~na614_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x71y97     80'h00_FE00_80_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a795_1 ( .OUT(na795_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7015_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a795_2 ( .OUT(na795_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na795_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a795_4 ( .OUT(na795_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na7014_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a795_5 ( .OUT(na795_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na795_2_i) );
// C_MX4b/D///      x92y78     80'h00_FE00_00_0040_0AC4_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_1 ( .OUT(na796_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na797_1),
                     .IN8(na796_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_2 ( .OUT(na796_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na796_1_i) );
// C_ORAND////      x78y73     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na155_1), .IN6(1'b0), .IN7(na354_2), .IN8(na9337_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x71y72     80'h00_0060_00_0000_0C08_FF31
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a798_4 ( .OUT(na798_2), .IN1(~na356_2), .IN2(~na5402_1), .IN3(1'b1), .IN4(~na5403_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x77y89     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a799_1 ( .OUT(na799_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na800_1), .IN8(na3914_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a799_5 ( .OUT(na799_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na799_1) );
// C_MX2b////      x70y77     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a800_1 ( .OUT(na800_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na5840_1), .IN8(na801_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x58y110     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a801_1 ( .OUT(na801_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2203_1), .IN7(1'b0), .IN8(~na624_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x81y91     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a803_1 ( .OUT(na803_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na804_1), .IN8(na3914_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a803_5 ( .OUT(na803_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na803_1) );
// C_MX2b////      x76y77     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a804_1 ( .OUT(na804_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na805_1), .IN8(~na3947_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y105     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a805_1 ( .OUT(na805_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2205_1), .IN7(1'b0), .IN8(~na1600_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x70y98     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a806_1 ( .OUT(na806_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7018_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a806_2 ( .OUT(na806_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na806_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a806_4 ( .OUT(na806_2_i), .IN1(1'b1), .IN2(na7017_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a806_5 ( .OUT(na806_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na806_2_i) );
// C_MX2b////D      x80y87     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a807_1 ( .OUT(na807_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3916_2), .IN8(~na808_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a807_5 ( .OUT(na807_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na807_1) );
// C_MX2b////      x70y104     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a808_1 ( .OUT(na808_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3949_1), .IN8(na809_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y108     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2209_1), .IN7(1'b0), .IN8(~na634_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x72y98     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a810_1 ( .OUT(na810_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7019_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a810_2 ( .OUT(na810_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na810_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a810_4 ( .OUT(na810_2_i), .IN1(na7234_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a810_5 ( .OUT(na810_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na810_2_i) );
// C_MX2b////D      x79y91     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a811_1 ( .OUT(na811_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na812_1), .IN8(na3918_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a811_5 ( .OUT(na811_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na811_1) );
// C_MX2b////      x72y107     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a812_1 ( .OUT(na812_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na5844_2), .IN8(na813_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x58y116     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a813_1 ( .OUT(na813_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2211_1), .IN7(1'b0), .IN8(~na1583_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x74y94     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a815_1 ( .OUT(na815_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3921_1), .IN8(~na816_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a815_5 ( .OUT(na815_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na815_1) );
// C_MX2b////      x72y106     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a816_1 ( .OUT(na816_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na5846_2), .IN6(na817_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x59y114     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2215_1), .IN7(1'b0), .IN8(~na664_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x77y91     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a819_1 ( .OUT(na819_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na820_1), .IN8(na3918_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a819_5 ( .OUT(na819_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na819_1) );
// C_MX2b////      x70y103     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a820_1 ( .OUT(na820_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na821_1), .IN8(~na3952_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y107     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a821_1 ( .OUT(na821_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2213_1), .IN7(1'b0), .IN8(~na658_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x73y98     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a822_1 ( .OUT(na822_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7022_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a822_2 ( .OUT(na822_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na822_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a822_4 ( .OUT(na822_2_i), .IN1(1'b1), .IN2(na7020_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a822_5 ( .OUT(na822_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na822_2_i) );
// C_MX2b////D      x72y96     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a823_1 ( .OUT(na823_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3921_2), .IN8(~na824_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a823_5 ( .OUT(na823_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na823_1) );
// C_MX2b////      x66y106     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a824_1 ( .OUT(na824_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3954_1), .IN8(na825_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x58y108     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a825_1 ( .OUT(na825_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2217_1), .IN7(1'b0), .IN8(~na669_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x74y99     80'h00_FE00_80_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a826_1 ( .OUT(na826_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na7023_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a826_2 ( .OUT(na826_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na826_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a826_4 ( .OUT(na826_2_i), .IN1(na7021_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a826_5 ( .OUT(na826_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na826_2_i) );
// C_MX4b/D///      x109y84     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9340_2),
                     .IN8(na3048_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_2 ( .OUT(na827_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na827_1_i) );
// C_MX2b////D      x76y95     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a828_1 ( .OUT(na828_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na829_1), .IN8(na3923_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a828_5 ( .OUT(na828_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na828_1) );
// C_MX2b////      x64y105     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a829_1 ( .OUT(na829_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na830_1), .IN8(~na3956_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x58y109     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a830_1 ( .OUT(na830_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2221_1), .IN7(1'b0), .IN8(~na679_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x68y98     80'h00_FE00_80_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a831_1 ( .OUT(na831_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na7024_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a831_2 ( .OUT(na831_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na831_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a831_4 ( .OUT(na831_2_i), .IN1(1'b1), .IN2(na7233_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a831_5 ( .OUT(na831_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na831_2_i) );
// C_MX4b/D///      x104y82     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a832_1 ( .OUT(na832_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na833_1),
                     .IN8(na832_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a832_2 ( .OUT(na832_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na832_1_i) );
// C_AND////      x104y85     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a833_1 ( .OUT(na833_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(na2532_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x74y96     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a834_1 ( .OUT(na834_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3925_1), .IN8(~na835_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a834_5 ( .OUT(na834_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na834_1) );
// C_MX2b////      x56y94     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a835_1 ( .OUT(na835_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na5850_2), .IN6(na836_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x59y120     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a836_1 ( .OUT(na836_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2223_1), .IN7(1'b0), .IN8(~na684_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x86y76     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a838_1 ( .OUT(na838_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2550_1),
                     .IN8(na838_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a838_2 ( .OUT(na838_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na838_1_i) );
// C_AND/D///      x106y86     80'h00_FE00_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_1 ( .OUT(na839_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na981_1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_2 ( .OUT(na839_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na839_1_i) );
// C_///AND/      x118y68     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a841_4 ( .OUT(na841_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na3219_2), .IN4(~na3227_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x77y94     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a843_1 ( .OUT(na843_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na844_1), .IN8(na3927_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a843_5 ( .OUT(na843_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na843_1) );
// C_MX2b////      x62y89     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a844_1 ( .OUT(na844_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na5852_1), .IN8(na845_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y118     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a845_1 ( .OUT(na845_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2227_1), .IN7(1'b0), .IN8(~na694_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x76y94     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_1 ( .OUT(na847_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3929_1), .IN8(~na848_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a847_5 ( .OUT(na847_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na847_1) );
// C_MX2b////      x72y110     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a848_1 ( .OUT(na848_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b0), .IN4(1'b0), .IN5(na849_1), .IN6(~na5854_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x61y117     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a849_1 ( .OUT(na849_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2231_1), .IN7(1'b0), .IN8(~na704_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x100y89     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a851_4 ( .OUT(na851_2_i), .IN1(na7029_1), .IN2(~na7028_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a851_5 ( .OUT(na851_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na851_2_i) );
// C_///AND/      x99y87     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a853_4 ( .OUT(na853_2), .IN1(na854_1), .IN2(1'b1), .IN3(na430_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y75     80'h00_0018_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a854_1 ( .OUT(na854_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na86_1), .IN6(na9154_2), .IN7(na8_1), .IN8(~na61_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y87     80'h00_0018_00_0000_0888_312F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a855_1 ( .OUT(na855_1), .IN1(1'b1), .IN2(1'b1), .IN3(na430_1), .IN4(~na452_2), .IN5(~na488_2), .IN6(~na435_1), .IN7(1'b1),
                     .IN8(~na452_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x100y80     80'h00_0060_00_0000_0C0E_FF5A
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a856_4 ( .OUT(na856_2), .IN1(na488_2), .IN2(1'b0), .IN3(~na430_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x79y90     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_1 ( .OUT(na857_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na858_1), .IN8(na3927_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a857_5 ( .OUT(na857_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na857_1) );
// C_MX2b////      x64y107     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a858_1 ( .OUT(na858_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na859_1), .IN8(~na3960_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y111     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a859_1 ( .OUT(na859_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2229_1), .IN7(1'b0), .IN8(~na699_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x69y101     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a860_1 ( .OUT(na860_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9216_2), .IN6(1'b1), .IN7(na7031_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a860_2 ( .OUT(na860_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na860_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a860_4 ( .OUT(na860_2_i), .IN1(na7026_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a860_5 ( .OUT(na860_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na860_2_i) );
// C_///ORAND/D      x96y92     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a861_4 ( .OUT(na861_2_i), .IN1(~na7032_1), .IN2(na7033_2), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a861_5 ( .OUT(na861_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na861_2_i) );
// C_MX2b////D      x78y96     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a863_1 ( .OUT(na863_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3929_2), .IN8(~na864_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a863_5 ( .OUT(na863_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na863_1) );
// C_MX2b////      x68y108     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a864_1 ( .OUT(na864_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3963_1), .IN8(na865_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y110     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a865_1 ( .OUT(na865_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2233_1), .IN7(1'b0), .IN8(~na719_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x68y99     80'h00_FE00_80_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a866_1 ( .OUT(na866_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na7034_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a866_2 ( .OUT(na866_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na866_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a866_4 ( .OUT(na866_2_i), .IN1(na7027_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a866_5 ( .OUT(na866_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na866_2_i) );
// C_MX4b/D///      x111y81     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a867_1 ( .OUT(na867_1_i), .IN1(1'b1), .IN2(na981_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na867_1), .IN6(na4177_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a867_2 ( .OUT(na867_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na867_1_i) );
// C_MX4b/D///      x113y81     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_1 ( .OUT(na868_1_i), .IN1(1'b1), .IN2(na981_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na868_1), .IN6(na4179_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_2 ( .OUT(na868_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na868_1_i) );
// C_MX4b/D///      x113y77     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1_i), .IN1(1'b1), .IN2(na981_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na869_1), .IN6(na4179_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_2 ( .OUT(na869_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na869_1_i) );
// C_ORAND/D//AND/D      x96y86     80'h00_FE00_80_0000_0C88_3E8F
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_1 ( .OUT(na870_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7036_1), .IN6(na871_2), .IN7(1'b0), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_2 ( .OUT(na870_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na870_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a870_4 ( .OUT(na870_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na904_1), .IN4(na870_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a870_5 ( .OUT(na870_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na870_2_i) );
// C_///ORAND/      x95y84     80'h00_0060_00_0000_0C08_FF7C
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a871_4 ( .OUT(na871_2), .IN1(1'b0), .IN2(na9347_2), .IN3(~na907_2), .IN4(~na872_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x102y82     80'h00_FE00_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a872_1 ( .OUT(na872_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na873_2), .IN7(na567_1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a872_2 ( .OUT(na872_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na872_1_i) );
// C_///AND/      x99y78     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a873_4 ( .OUT(na873_2), .IN1(1'b1), .IN2(na874_1), .IN3(na436_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y80     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a874_1 ( .OUT(na874_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na566_1), .IN6(na435_2), .IN7(1'b1), .IN8(na9228_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y81     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_1 ( .OUT(na875_1_i), .IN1(na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na875_1),
                     .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_2 ( .OUT(na875_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na875_1_i) );
// C_AND////      x99y77     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a876_1 ( .OUT(na876_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(na873_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x105y79     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_1 ( .OUT(na877_1_i), .IN1(na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na877_1), .IN6(na259_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_2 ( .OUT(na877_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na877_1_i) );
// C_AND/D//AND/D      x73y83     80'h00_FA00_80_0000_0C88_F8CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_1 ( .OUT(na878_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na878_2), .IN6(na410_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_2 ( .OUT(na878_1), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na878_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a878_4 ( .OUT(na878_2_i), .IN1(1'b1), .IN2(na410_1), .IN3(1'b1), .IN4(na984_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a878_5 ( .OUT(na878_2), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na878_2_i) );
// C_MX4b/D///      x107y77     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a879_1 ( .OUT(na879_1_i), .IN1(na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na879_1), .IN6(na262_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a879_2 ( .OUT(na879_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na879_1_i) );
// C_MX4b/D///      x98y76     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a880_1 ( .OUT(na880_1_i), .IN1(~na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                     .IN8(na880_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a880_2 ( .OUT(na880_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na880_1_i) );
// C_MX4b/D///      x112y82     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a881_1 ( .OUT(na881_1_i), .IN1(~na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                     .IN8(na881_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a881_2 ( .OUT(na881_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na881_1_i) );
// C_MX4b/D///      x111y77     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a882_1 ( .OUT(na882_1_i), .IN1(na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na882_1), .IN6(na265_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a882_2 ( .OUT(na882_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na882_1_i) );
// C_MX4b/D///      x110y84     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_1 ( .OUT(na883_1_i), .IN1(1'b1), .IN2(~na981_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na4175_1),
                     .IN8(na883_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_2 ( .OUT(na883_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na883_1_i) );
// C_ORAND/D///      x98y88     80'h00_FE00_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a884_1 ( .OUT(na884_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7038_2), .IN6(na7039_1), .IN7(na855_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a884_2 ( .OUT(na884_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na884_1_i) );
// C_ORAND/D///      x99y96     80'h00_FE00_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a886_1 ( .OUT(na886_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7041_1), .IN6(~na7040_2), .IN7(na855_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a886_2 ( .OUT(na886_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na886_1_i) );
// C_///ORAND/D      x102y91     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a888_4 ( .OUT(na888_2_i), .IN1(na7043_2), .IN2(~na7042_2), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a888_5 ( .OUT(na888_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na888_2_i) );
// C_MX4b/D///      x101y94     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a890_1 ( .OUT(na890_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na581_1), .IN6(na890_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a890_2 ( .OUT(na890_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na890_1_i) );
// C_MX4b/D///      x105y75     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1_i), .IN1(1'b1), .IN2(na161_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na891_1), .IN6(na6477_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_2 ( .OUT(na891_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na891_1_i) );
// C_MX4b/D///      x105y84     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a892_1 ( .OUT(na892_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9349_2), .IN6(na893_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a892_2 ( .OUT(na892_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na892_1_i) );
// C_///AND/      x109y78     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a893_4 ( .OUT(na893_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1113_1), .IN4(na2528_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x100y92     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a894_1 ( .OUT(na894_1_i), .IN1(~na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                     .IN8(na894_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a894_2 ( .OUT(na894_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na894_1_i) );
// C_MX4b/D///      x93y87     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a895_1 ( .OUT(na895_1_i), .IN1(na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na895_1), .IN6(na265_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a895_2 ( .OUT(na895_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na895_1_i) );
// C_AND/D///      x100y96     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a896_1 ( .OUT(na896_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1860_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a896_2 ( .OUT(na896_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na896_1_i) );
// C_MX4b/D///      x100y90     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1_i), .IN1(~na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                     .IN8(na897_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_2 ( .OUT(na897_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na897_1_i) );
// C_AND////      x115y77     80'h00_0018_00_0000_0888_4554
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a898_1 ( .OUT(na898_1), .IN1(~na3256_1), .IN2(na3345_1), .IN3(~na9810_2), .IN4(1'b1), .IN5(~na3352_2), .IN6(1'b1), .IN7(~na3596_2),
                     .IN8(na3590_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x121y71     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_1 ( .OUT(na900_1_i), .IN1(na898_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na900_1), .IN6(na901_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a900_2 ( .OUT(na900_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na900_1_i) );
// C_AND////      x123y70     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a901_1 ( .OUT(na901_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na900_1), .IN6(na7044_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x97y89     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a902_1 ( .OUT(na902_1_i), .IN1(na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na902_1), .IN6(na262_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a902_2 ( .OUT(na902_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na902_1_i) );
// C_MX4b/D///      x90y75     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a903_1 ( .OUT(na903_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na903_1),
                     .IN8(na2548_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a903_2 ( .OUT(na903_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na903_1_i) );
// C_AND/D///      x98y83     80'h00_FE00_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a904_1 ( .OUT(na904_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na905_1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a904_2 ( .OUT(na904_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na904_1_i) );
// C_MX2a////      x102y89     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a905_1 ( .OUT(na905_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na904_1), .IN4(~na159_1), .IN5(na906_1), .IN6(na873_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y75     80'h00_0018_00_0000_0C88_82FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a906_1 ( .OUT(na906_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na854_1), .IN6(~na36_1), .IN7(na489_1), .IN8(na9948_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x106y81     80'h00_FE00_80_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a907_4 ( .OUT(na907_2_i), .IN1(1'b1), .IN2(~na908_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a907_5 ( .OUT(na907_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na907_2_i) );
// C_MX2a////      x95y86     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a908_1 ( .OUT(na908_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na907_2), .IN4(~na159_1), .IN5(na9266_2), .IN6(na873_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x89y96     80'h00_FE00_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a909_1 ( .OUT(na909_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7046_1), .IN6(na7047_1), .IN7(na855_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a909_2 ( .OUT(na909_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na909_1_i) );
// C_///AND/D      x111y88     80'h00_FE00_80_0000_0C08_FF38
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a911_4 ( .OUT(na911_2_i), .IN1(na853_2), .IN2(na873_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a911_5 ( .OUT(na911_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na911_2_i) );
// C_MX4b/D///      x107y75     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a912_1 ( .OUT(na912_1_i), .IN1(1'b1), .IN2(na981_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na912_1), .IN6(na4173_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a912_2 ( .OUT(na912_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na912_1_i) );
// C_AND/D//AND/D      x90y93     80'h00_FE00_80_0000_0C88_351F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a913_1 ( .OUT(na913_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na914_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a913_2 ( .OUT(na913_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na913_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a913_4 ( .OUT(na913_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1875_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a913_5 ( .OUT(na913_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na913_2_i) );
// C_MX2a////      x89y83     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a914_1 ( .OUT(na914_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na913_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na915_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y86     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a915_4 ( .OUT(na915_2), .IN1(na9954_2), .IN2(na435_1), .IN3(na436_1), .IN4(~na452_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x89y80     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a916_1 ( .OUT(na916_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9355_2),
                     .IN8(na2547_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a916_2 ( .OUT(na916_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na916_1_i) );
// C_MX4b/D///      x87y71     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a917_1 ( .OUT(na917_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na917_1), .IN6(na2546_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a917_2 ( .OUT(na917_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na917_1_i) );
// C_MX4b/D///      x87y77     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a918_1 ( .OUT(na918_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na918_1), .IN6(na2545_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a918_2 ( .OUT(na918_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na918_1_i) );
// C_MX4b/D///      x89y77     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a919_1 ( .OUT(na919_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na919_1), .IN6(na2544_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a919_2 ( .OUT(na919_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na919_1_i) );
// C_MX4b/D///      x88y75     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_1 ( .OUT(na920_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na920_1),
                     .IN8(na2543_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_2 ( .OUT(na920_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na920_1_i) );
// C_MX4b/D///      x92y76     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a921_1 ( .OUT(na921_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2542_1),
                     .IN8(na921_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a921_2 ( .OUT(na921_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na921_1_i) );
// C_MX2a////      x87y88     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a923_1 ( .OUT(na923_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na925_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na924_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y86     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a924_1 ( .OUT(na924_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9954_2), .IN6(na435_1), .IN7(na433_2), .IN8(na9230_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x94y93     80'h00_FE00_80_0000_0C88_1F33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a925_1 ( .OUT(na925_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na926_1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a925_2 ( .OUT(na925_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na925_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a925_4 ( .OUT(na925_2_i), .IN1(1'b1), .IN2(~na923_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a925_5 ( .OUT(na925_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na925_2_i) );
// C_MX2a////      x116y97     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a926_1 ( .OUT(na926_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na925_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na924_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x95y94     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a927_4 ( .OUT(na927_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na928_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a927_5 ( .OUT(na927_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na927_2_i) );
// C_MX2a////      x88y99     80'h00_0018_00_0040_0CAA_8F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a928_1 ( .OUT(na928_1), .IN1(1'b0), .IN2(~na927_2), .IN3(1'b0), .IN4(~na159_1), .IN5(1'b1), .IN6(1'b1), .IN7(na436_1), .IN8(na929_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y84     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a929_4 ( .OUT(na929_2), .IN1(na9954_2), .IN2(na435_1), .IN3(na433_1), .IN4(na9223_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x98y93     80'h00_FE00_00_0040_0AC3_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a930_1 ( .OUT(na930_1_i), .IN1(na931_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na930_1),
                     .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a930_2 ( .OUT(na930_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na930_1_i) );
// C_AND////      x93y91     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a931_1 ( .OUT(na931_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na488_1), .IN6(na932_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y88     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a932_1 ( .OUT(na932_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(~na435_1), .IN7(na436_1), .IN8(~na452_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y89     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a933_1 ( .OUT(na933_1_i), .IN1(na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na933_1),
                     .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a933_2 ( .OUT(na933_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na933_1_i) );
// C_///AND/      x103y83     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a934_4 ( .OUT(na934_2), .IN1(na428_1), .IN2(na932_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y89     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a935_1 ( .OUT(na935_1_i), .IN1(na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na935_1), .IN6(na259_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a935_2 ( .OUT(na935_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na935_1_i) );
// C_MX4b/D///      x101y93     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a936_1 ( .OUT(na936_1_i), .IN1(~na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                     .IN8(na9358_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a936_2 ( .OUT(na936_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na936_1_i) );
// C_MX4b/D///      x102y92     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a937_1 ( .OUT(na937_1_i), .IN1(~na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                     .IN8(na937_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a937_2 ( .OUT(na937_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na937_1_i) );
// C_MX4b/D///      x103y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a938_1 ( .OUT(na938_1_i), .IN1(na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na938_1), .IN6(na262_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a938_2 ( .OUT(na938_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na938_1_i) );
// C_MX4b/D///      x104y90     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a939_1 ( .OUT(na939_1_i), .IN1(~na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                     .IN8(na939_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a939_2 ( .OUT(na939_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na939_1_i) );
// C_MX4b/D///      x110y94     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a940_1 ( .OUT(na940_1_i), .IN1(~na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                     .IN8(na940_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a940_2 ( .OUT(na940_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na940_1_i) );
// C_MX4b/D///      x93y93     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a941_1 ( .OUT(na941_1_i), .IN1(na934_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na941_1), .IN6(na265_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a941_2 ( .OUT(na941_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na941_1_i) );
// C_AND/D///      x93y62     80'h00_FE00_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a942_1 ( .OUT(na942_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na943_1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a942_2 ( .OUT(na942_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na942_1_i) );
// C_MX2a////      x91y80     80'h00_0018_00_0040_0CAA_8F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a943_1 ( .OUT(na943_1), .IN1(1'b0), .IN2(~na942_1), .IN3(1'b0), .IN4(~na159_1), .IN5(1'b1), .IN6(1'b1), .IN7(na436_1), .IN8(na944_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y78     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a944_1 ( .OUT(na944_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(na435_1), .IN7(na9222_2), .IN8(~na452_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x116y69     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_1 ( .OUT(na945_1_i), .IN1(na946_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na945_1),
                     .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_2 ( .OUT(na945_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na945_1_i) );
// C_///AND/      x111y69     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a946_4 ( .OUT(na946_2), .IN1(1'b1), .IN2(1'b1), .IN3(na436_1), .IN4(na947_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y76     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a947_1 ( .OUT(na947_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(na435_1), .IN7(na433_1), .IN8(na9223_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x119y67     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a948_1 ( .OUT(na948_1_i), .IN1(na946_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na948_1), .IN6(na259_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a948_2 ( .OUT(na948_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na948_1_i) );
// C_MX4b/D///      x118y70     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a949_1 ( .OUT(na949_1_i), .IN1(~na946_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                     .IN8(na949_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a949_2 ( .OUT(na949_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na949_1_i) );
// C_AND/D//AND/D      x118y104     80'h00_FE00_80_0000_0C88_CACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a950_1 ( .OUT(na950_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6486_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a950_2 ( .OUT(na950_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na950_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a950_4 ( .OUT(na950_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na950_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a950_5 ( .OUT(na950_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na950_2_i) );
// C_AND///AND/      x119y99     80'h00_0078_00_0000_0C88_3281
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a951_1 ( .OUT(na951_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2987_1), .IN6(~na2983_1), .IN7(1'b1), .IN8(~na238_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a951_4 ( .OUT(na951_2), .IN1(~na1010_1), .IN2(~na9377_2), .IN3(na1013_1), .IN4(na1018_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x116y104     80'h00_FE00_80_0000_0C88_F8CF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a952_1 ( .OUT(na952_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(na6487_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a952_2 ( .OUT(na952_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na952_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a952_4 ( .OUT(na952_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na952_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a952_5 ( .OUT(na952_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na952_2_i) );
// C_AND/D///      x108y93     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a953_1 ( .OUT(na953_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na954_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a953_2 ( .OUT(na953_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na953_1_i) );
// C_AND////      x107y91     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a954_1 ( .OUT(na954_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na932_1), .IN7(1'b1), .IN8(na9362_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y78     80'h00_0018_00_0000_0888_A4C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a955_1 ( .OUT(na955_1), .IN1(1'b1), .IN2(~na431_1), .IN3(1'b1), .IN4(na6673_2), .IN5(~na86_1), .IN6(na36_2), .IN7(na489_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x117y103     80'h00_FE00_80_0000_0C88_AAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a957_1 ( .OUT(na957_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(na6488_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a957_2 ( .OUT(na957_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na957_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a957_4 ( .OUT(na957_2_i), .IN1(na957_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a957_5 ( .OUT(na957_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na957_2_i) );
// C_MX4b/D///      x117y68     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a958_1 ( .OUT(na958_1_i), .IN1(~na946_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                     .IN8(na9363_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a958_2 ( .OUT(na958_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na958_1_i) );
// C_AND/D//AND/D      x114y104     80'h00_FE00_80_0000_0C88_F8CF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a959_1 ( .OUT(na959_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(na6489_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a959_2 ( .OUT(na959_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na959_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a959_4 ( .OUT(na959_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na959_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a959_5 ( .OUT(na959_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na959_2_i) );
// C_MX4b/D///      x97y99     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a960_1 ( .OUT(na960_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na960_1), .IN6(na961_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a960_2 ( .OUT(na960_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na960_1_i) );
// C_///AND/      x89y82     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a961_4 ( .OUT(na961_2), .IN1(na2540_1), .IN2(1'b1), .IN3(~na1113_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x89y74     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a962_1 ( .OUT(na962_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2541_1), .IN6(na962_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a962_2 ( .OUT(na962_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na962_1_i) );
// C_MX4b/D///      x90y78     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a963_1 ( .OUT(na963_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2539_1),
                     .IN8(na963_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a963_2 ( .OUT(na963_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na963_1_i) );
// C_AND/D//AND/D      x116y103     80'h00_FE00_80_0000_0C88_CAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a964_1 ( .OUT(na964_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6490_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a964_2 ( .OUT(na964_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na964_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a964_4 ( .OUT(na964_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na964_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a964_5 ( .OUT(na964_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na964_2_i) );
// C_AND/D//AND/D      x122y103     80'h00_FE00_80_0000_0C88_F8AF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a965_1 ( .OUT(na965_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(na6491_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a965_2 ( .OUT(na965_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na965_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a965_4 ( .OUT(na965_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na965_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a965_5 ( .OUT(na965_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na965_2_i) );
// C_AND/D//AND/D      x116y106     80'h00_FE00_80_0000_0C88_AACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a966_1 ( .OUT(na966_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(na6492_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a966_2 ( .OUT(na966_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na966_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a966_4 ( .OUT(na966_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na966_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a966_5 ( .OUT(na966_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na966_2_i) );
// C_AND/D//AND/D      x118y107     80'h00_FE00_80_0000_0C88_CAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a967_1 ( .OUT(na967_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6493_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a967_2 ( .OUT(na967_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na967_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a967_4 ( .OUT(na967_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na967_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a967_5 ( .OUT(na967_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na967_2_i) );
// C_AND/D//AND/D      x119y103     80'h00_FE00_80_0000_0C88_AAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a968_1 ( .OUT(na968_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(na6494_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a968_2 ( .OUT(na968_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na968_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a968_4 ( .OUT(na968_2_i), .IN1(na968_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a968_5 ( .OUT(na968_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na968_2_i) );
// C_AND/D//AND/D      x114y103     80'h00_FE00_80_0000_0C88_CAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a969_1 ( .OUT(na969_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6495_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a969_2 ( .OUT(na969_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na969_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a969_4 ( .OUT(na969_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na969_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a969_5 ( .OUT(na969_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na969_2_i) );
// C_AND/D//AND/D      x113y103     80'h00_FE00_80_0000_0C88_AAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a970_1 ( .OUT(na970_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na951_1), .IN6(1'b1), .IN7(na6496_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a970_2 ( .OUT(na970_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na970_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a970_4 ( .OUT(na970_2_i), .IN1(na970_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a970_5 ( .OUT(na970_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na970_2_i) );
// C_ORAND/D///      x53y111     80'h00_FE00_00_0000_0888_3F5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a971_1 ( .OUT(na971_1_i), .IN1(na971_1), .IN2(na7049_2), .IN3(~na409_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(~na6626_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a971_2 ( .OUT(na971_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na971_1_i) );
// C_ORAND/D///      x118y48     80'h00_FE00_00_0000_0888_EF33
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_1 ( .OUT(na973_1_i), .IN1(1'b0), .IN2(~na974_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na9730_2),
                     .IN8(na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_2 ( .OUT(na973_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na973_1_i) );
// C_AND////      x117y52     80'h00_0018_00_0000_0888_238C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a974_1 ( .OUT(na974_1), .IN1(1'b1), .IN2(na3031_2), .IN3(na9364_2), .IN4(na3032_2), .IN5(1'b1), .IN6(~na3031_1), .IN7(na1223_1),
                     .IN8(~na3032_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x84y65     80'h00_FE00_80_0000_0C88_3C28
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a977_1 ( .OUT(na977_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na467_1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a977_2 ( .OUT(na977_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na977_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a977_4 ( .OUT(na977_2_i), .IN1(na468_1), .IN2(na27_1), .IN3(na469_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a977_5 ( .OUT(na977_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na977_2_i) );
// C_AND/D///      x90y69     80'h00_FE00_00_0000_0888_3C2C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a978_1 ( .OUT(na978_1_i), .IN1(1'b1), .IN2(na18_1), .IN3(na469_1), .IN4(~na28_1), .IN5(1'b1), .IN6(na27_1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a978_2 ( .OUT(na978_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na978_1_i) );
// C_AND/D///      x97y76     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a979_1 ( .OUT(na979_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a979_2 ( .OUT(na979_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na979_1_i) );
// C_MX4b/D///      x113y98     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a980_1 ( .OUT(na980_1_i), .IN1(~na951_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na7051_1), .IN6(na980_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a980_2 ( .OUT(na980_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na980_1_i) );
// C_AND/D///      x111y82     80'h00_FE00_00_0000_0888_8514
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a981_1 ( .OUT(na981_1_i), .IN1(~na3256_1), .IN2(na3345_1), .IN3(~na4204_2), .IN4(~na6626_1), .IN5(~na3290_1), .IN6(1'b1),
                     .IN7(na3596_2), .IN8(na983_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a981_2 ( .OUT(na981_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na981_1_i) );
// C_AND////      x116y74     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a983_1 ( .OUT(na983_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3352_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na3590_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x76y82     80'h00_FA00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a984_1 ( .OUT(na984_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na410_1), .IN7(1'b1), .IN8(na984_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a984_2 ( .OUT(na984_1), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na984_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a984_4 ( .OUT(na984_2_i), .IN1(1'b1), .IN2(na410_1), .IN3(1'b1), .IN4(na999_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a984_5 ( .OUT(na984_2), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na984_2_i) );
// C_AND/D//AND/D      x125y49     80'h00_FE00_80_0000_0C88_1F55
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a985_1 ( .OUT(na985_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na986_1), .IN8(~na988_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a985_2 ( .OUT(na985_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na985_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a985_4 ( .OUT(na985_2_i), .IN1(~na2800_1), .IN2(1'b1), .IN3(~na986_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a985_5 ( .OUT(na985_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na985_2_i) );
// C_AND////      x122y61     80'h00_0018_00_0000_0888_4351
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a986_1 ( .OUT(na986_1), .IN1(~na3594_1), .IN2(~na3356_1), .IN3(~na3219_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na3222_1), .IN7(~na3219_1),
                     .IN8(na3227_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x130y50     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a988_1 ( .OUT(na988_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na500_2), .IN5(~na985_1), .IN6(1'b0), .IN7(~na7052_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y48     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a989_1 ( .OUT(na989_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na985_1), .IN6(na2972_2), .IN7(na9371_2), .IN8(na9725_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x111y89     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a990_1 ( .OUT(na990_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na990_1), .IN6(na991_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a990_2 ( .OUT(na990_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na990_1_i) );
// C_///AND/      x103y80     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a991_4 ( .OUT(na991_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1113_1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y95     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a992_1 ( .OUT(na992_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na992_1), .IN6(na993_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a992_2 ( .OUT(na992_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na992_1_i) );
// C_AND////      x93y84     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a993_1 ( .OUT(na993_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2541_1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x119y95     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_1 ( .OUT(na995_1_i), .IN1(1'b1), .IN2(na996_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na995_1), .IN6(~na998_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_2 ( .OUT(na995_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na995_1_i) );
// C_///ANDXOR/      x117y96     80'h00_0060_00_0000_0C06_FF57
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a996_4 ( .OUT(na996_2), .IN1(na951_1), .IN2(na1064_1), .IN3(na997_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x112y91     80'h00_0018_00_0040_0C55_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a997_1 ( .OUT(na997_1), .IN1(~na7054_1), .IN2(1'b0), .IN3(~na7055_1), .IN4(1'b0), .IN5(na7054_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na9703_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x119y96     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a998_1 ( .OUT(na998_1), .IN1(1'b0), .IN2(1'b0), .IN3(na997_1), .IN4(1'b1), .IN5(~na3972_2), .IN6(1'b0), .IN7(~na3865_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x74y82     80'h00_FA00_80_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_1 ( .OUT(na999_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na410_1), .IN7(1'b1), .IN8(na999_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_2 ( .OUT(na999_1), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na999_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a999_4 ( .OUT(na999_2_i), .IN1(1'b1), .IN2(na410_1), .IN3(na4853_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a999_5 ( .OUT(na999_2), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na999_2_i) );
// C_MX4b/D///      x88y80     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2538_1),
                      .IN8(na1000_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_2 ( .OUT(na1000_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1000_1_i) );
// C_MX4b/D///      x84y76     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1001_1 ( .OUT(na1001_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2537_1), .IN6(na9375_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1001_2 ( .OUT(na1001_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1001_1_i) );
// C_MX4b/D///      x86y77     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1002_1 ( .OUT(na1002_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1002_1),
                      .IN8(na2536_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1002_2 ( .OUT(na1002_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1002_1_i) );
// C_MX4b/D///      x92y80     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_1 ( .OUT(na1003_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2534_2),
                      .IN8(na1003_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_2 ( .OUT(na1003_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1003_1_i) );
// C_MX4b/D///      x90y77     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1004_1 ( .OUT(na1004_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1004_1),
                      .IN8(na2532_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1004_2 ( .OUT(na1004_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1004_1_i) );
// C_MX4b/D///      x90y79     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1005_1 ( .OUT(na1005_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1005_1),
                      .IN8(na2530_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1005_2 ( .OUT(na1005_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1005_1_i) );
// C_///ICOMP/D      x111y87     80'h00_FE00_80_0000_0C08_FF36
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1006_4 ( .OUT(na1006_2_i), .IN1(na1006_2), .IN2(~na9374_2), .IN3(1'b0), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1006_5 ( .OUT(na1006_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1006_2_i) );
// C_MX4b/D///      x111y92     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1007_1 ( .OUT(na1007_1_i), .IN1(~na9373_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na7057_2), .IN6(na1007_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1007_2 ( .OUT(na1007_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1007_1_i) );
// C_///ICOMP/D      x105y80     80'h00_FE00_80_0000_0C08_FF39
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1008_4 ( .OUT(na1008_2_i), .IN1(~na10027_2), .IN2(~na1008_2), .IN3(1'b0), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1008_5 ( .OUT(na1008_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1008_2_i) );
// C_MX4b/D///      x108y76     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1_i), .IN1(na10027_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na7059_1),
                      .IN8(na1009_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_2 ( .OUT(na1009_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1009_1_i) );
// C_MX4b/D///      x121y83     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_1 ( .OUT(na1010_1_i), .IN1(na1011_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1010_1), .IN6(~na9376_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_2 ( .OUT(na1010_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1010_1_i) );
// C_///XOR/      x119y81     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1011_4 ( .OUT(na1011_2), .IN1(na10027_2), .IN2(~na1012_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x119y78     80'h00_0018_00_0000_0C88_E5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_1 ( .OUT(na1012_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1014_2), .IN6(1'b0), .IN7(na1013_1), .IN8(na237_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x116y87     80'h00_FA18_00_0000_0888_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1013_1 ( .OUT(na1013_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2987_1), .IN6(na2983_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1013_5 ( .OUT(na1013_2), .CLK(na4116_1), .EN(na3339_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1013_1) );
// C_///AND/      x121y81     80'h00_0060_00_0000_0C08_FF45
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1014_4 ( .OUT(na1014_2), .IN1(~na1010_1), .IN2(1'b1), .IN3(~na1016_1), .IN4(na1018_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x122y81     80'h00_FE00_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_1 ( .OUT(na1016_1_i), .IN1(na1011_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1016_1),
                      .IN8(~na1017_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_2 ( .OUT(na1016_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1016_1_i) );
// C_MX2b////      x128y80     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1017_1 ( .OUT(na1017_1), .IN1(1'b1), .IN2(~na1012_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3868_1), .IN6(~na9860_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x122y82     80'h00_FE00_00_0040_0AC4_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_1 ( .OUT(na1018_1_i), .IN1(~na1011_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1019_1),
                      .IN8(na1018_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_2 ( .OUT(na1018_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1018_1_i) );
// C_MX2b////      x130y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1019_1 ( .OUT(na1019_1), .IN1(1'b1), .IN2(~na1012_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3868_2), .IN6(~na9861_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP/D///      x111y73     80'h00_FE00_00_0000_0C88_36FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1020_1 ( .OUT(na1020_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1020_1), .IN6(~na1012_1), .IN7(1'b0), .IN8(na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1020_2 ( .OUT(na1020_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1020_1_i) );
// C_MX4b/D///      x114y75     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1021_1 ( .OUT(na1021_1_i), .IN1(1'b1), .IN2(na1012_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1021_1),
                      .IN8(na7062_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1021_2 ( .OUT(na1021_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1021_1_i) );
// C_AND/D///      x105y95     80'h00_FE00_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_1 ( .OUT(na1022_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1023_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_2 ( .OUT(na1022_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1022_1_i) );
// C_MX2a////      x118y101     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_1 ( .OUT(na1023_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na9378_2), .IN4(~na159_1), .IN5(na853_2), .IN6(na1024_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y90     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1024_1 ( .OUT(na1024_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na566_1), .IN6(na435_1), .IN7(na436_1), .IN8(~na452_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x102y75     80'h00_FE00_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1026_1 ( .OUT(na1026_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1027_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1026_2 ( .OUT(na1026_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1026_1_i) );
// C_MX2a////      x102y73     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1027_1 ( .OUT(na1027_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1026_1), .IN4(~na159_1), .IN5(na1028_1), .IN6(na1024_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y75     80'h00_0018_00_0000_0888_A4C2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1), .IN1(na9947_2), .IN2(~na36_1), .IN3(1'b1), .IN4(na6673_2), .IN5(~na86_1), .IN6(na36_2), .IN7(na489_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x100y87     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1030_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_2 ( .OUT(na1030_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1030_1_i) );
// C_MX4b/D///      x101y91     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1032_1 ( .OUT(na1032_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1032_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1032_2 ( .OUT(na1032_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1032_1_i) );
// C_MX4b/D///      x116y107     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1_i), .IN1(1'b1), .IN2(~na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na9379_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_2 ( .OUT(na1033_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1033_1_i) );
// C_AND///AND/      x105y91     80'h00_0078_00_0000_0C88_5AAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1034_1 ( .OUT(na1034_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2522_1), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1034_4 ( .OUT(na1034_2), .IN1(1'b1), .IN2(na1024_1), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x113y107     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_1 ( .OUT(na1035_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na9380_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_2 ( .OUT(na1035_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1035_1_i) );
// C_///AND/D      x110y82     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1036_4 ( .OUT(na1036_2_i), .IN1(na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1036_5 ( .OUT(na1036_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1036_2_i) );
// C_///AND/      x111y85     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1037_4 ( .OUT(na1037_2), .IN1(na853_2), .IN2(1'b1), .IN3(na490_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x73y79     80'h00_FA00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1038_1 ( .OUT(na1038_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1038_2), .IN6(na410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1038_2 ( .OUT(na1038_1), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1038_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1038_4 ( .OUT(na1038_2_i), .IN1(na878_1), .IN2(na410_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1038_5 ( .OUT(na1038_2), .CLK(na4116_1), .EN(na410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1038_2_i) );
// C_MX4b/D///      x111y91     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1_i), .IN1(na954_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9381_2),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_2 ( .OUT(na1039_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1039_1_i) );
// C_AND/D///      x95y87     80'h00_FE00_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1040_1 ( .OUT(na1040_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9226_2), .IN6(~na7063_1), .IN7(na433_2),
                      .IN8(~na452_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1040_2 ( .OUT(na1040_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1040_1_i) );
// C_ORAND////      x107y86     80'h00_0018_00_0000_0888_3FAB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1042_1 ( .OUT(na1042_1), .IN1(na6828_1), .IN2(~na1525_2), .IN3(na9382_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(~na1046_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x87y73     80'h00_0060_00_0000_0C0E_FF0B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1045_4 ( .OUT(na1045_2), .IN1(na7068_1), .IN2(~na1525_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x88y74     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1046_4 ( .OUT(na1046_2), .IN1(1'b0), .IN2(na1525_2), .IN3(na63_1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x108y82     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1048_4 ( .OUT(na1048_2_i), .IN1(na1049_1), .IN2(na7071_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1048_5 ( .OUT(na1048_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1048_2_i) );
// C_AND////      x109y83     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1049_1 ( .OUT(na1049_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2926_1), .IN6(1'b1), .IN7(na298_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x109y68     80'h00_FE00_80_0000_0C88_4F3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1053_1 ( .OUT(na1053_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7076_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1053_2 ( .OUT(na1053_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1053_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1053_4 ( .OUT(na1053_2_i), .IN1(1'b1), .IN2(na1598_1), .IN3(1'b1), .IN4(~na7354_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1053_5 ( .OUT(na1053_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1053_2_i) );
// C_///AND/      x102y80     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1054_4 ( .OUT(na1054_2), .IN1(na7078_1), .IN2(na435_2), .IN3(na9224_2), .IN4(na9228_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y66     80'h00_0018_00_0000_0888_D355
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_1 ( .OUT(na1055_1), .IN1(~na488_1), .IN2(1'b0), .IN3(~na567_1), .IN4(1'b0), .IN5(1'b0), .IN6(~na955_1), .IN7(~na430_1),
                      .IN8(na9243_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x100y75     80'h00_FE00_80_0000_0C88_4FC8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1057_1 ( .OUT(na1057_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7082_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1057_2 ( .OUT(na1057_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1057_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1057_4 ( .OUT(na1057_2_i), .IN1(na428_1), .IN2(na1598_1), .IN3(1'b1), .IN4(na9122_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1057_5 ( .OUT(na1057_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1057_2_i) );
// C_AND/D//AND/D      x108y75     80'h00_FE00_80_0000_0C88_4FCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_1 ( .OUT(na1059_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7086_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_2 ( .OUT(na1059_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1059_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1059_4 ( .OUT(na1059_2_i), .IN1(1'b1), .IN2(na958_1), .IN3(1'b1), .IN4(na947_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1059_5 ( .OUT(na1059_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1059_2_i) );
// C_AND/D//AND/D      x98y95     80'h00_FE00_80_0000_0C88_351F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_1 ( .OUT(na1061_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1062_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_2 ( .OUT(na1061_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1061_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1061_4 ( .OUT(na1061_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1879_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1061_5 ( .OUT(na1061_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1061_2_i) );
// C_MX2a////      x95y95     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1062_1 ( .OUT(na1062_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1061_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1063_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y88     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_1 ( .OUT(na1063_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(na435_2), .IN7(na436_1), .IN8(~na9228_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//ICOMP/D      x115y96     80'h00_FE00_80_0000_0C88_3336
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1064_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_2 ( .OUT(na1064_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1064_1_i) );
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1064_4 ( .OUT(na1064_2_i), .IN1(~na9388_2), .IN2(na1064_1), .IN3(1'b0), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1064_5 ( .OUT(na1064_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1064_2_i) );
// C_AND/D//AND/D      x76y71     80'h00_FE00_80_0000_0C88_351F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1065_1 ( .OUT(na1065_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1066_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1065_2 ( .OUT(na1065_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1065_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1065_4 ( .OUT(na1065_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1872_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1065_5 ( .OUT(na1065_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1065_2_i) );
// C_MX2a////      x71y73     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1066_1 ( .OUT(na1066_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1065_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1067_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y84     80'h00_0060_00_0000_0C08_FF22
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1067_4 ( .OUT(na1067_2), .IN1(na566_1), .IN2(~na435_1), .IN3(na436_1), .IN4(~na452_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y105     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1068_1 ( .OUT(na1068_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1068_1), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1068_2 ( .OUT(na1068_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1068_1_i) );
// C_MX4b/D///      x111y107     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_1 ( .OUT(na1069_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na9392_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_2 ( .OUT(na1069_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1069_1_i) );
// C_MX4b/D///      x111y109     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na9393_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_2 ( .OUT(na1070_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1070_1_i) );
// C_MX4b/D///      x111y111     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_1 ( .OUT(na1071_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1071_1), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_2 ( .OUT(na1071_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1071_1_i) );
// C_MX4b/D///      x103y97     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1072_1 ( .OUT(na1072_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1072_1), .IN6(na1073_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1072_2 ( .OUT(na1072_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1072_1_i) );
// C_AND///AND/      x107y112     80'h00_0078_00_0000_0C88_5AF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1073_1 ( .OUT(na1073_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(~na1113_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1073_4 ( .OUT(na1073_2), .IN1(na428_1), .IN2(na1024_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x107y90     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1074_1 ( .OUT(na1074_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na1074_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1074_2 ( .OUT(na1074_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1074_1_i) );
// C_MX4b/D///      x99y93     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1075_1 ( .OUT(na1075_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1075_1), .IN6(na454_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1075_2 ( .OUT(na1075_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1075_1_i) );
// C_MX4b/D///      x87y81     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1076_1 ( .OUT(na1076_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1076_1), .IN6(na2524_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1076_2 ( .OUT(na1076_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1076_1_i) );
// C_MX4b/D///      x107y97     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1077_1 ( .OUT(na1077_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1077_1), .IN6(na1078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1077_2 ( .OUT(na1077_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1077_1_i) );
// C_AND////      x95y90     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1078_1 ( .OUT(na1078_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(na2526_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x118y102     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_1 ( .OUT(na1079_1_i), .IN1(1'b1), .IN2(~na454_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na833_1),
                      .IN8(na1079_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_2 ( .OUT(na1079_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1079_1_i) );
// C_MX4b/D///      x111y95     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1080_1 ( .OUT(na1080_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1080_1), .IN6(na893_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1080_2 ( .OUT(na1080_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1080_1_i) );
// C_MX4b/D///      x107y93     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na833_1),
                      .IN8(na9397_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_2 ( .OUT(na1081_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1081_1_i) );
// C_MX4b/D///      x87y80     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1082_1 ( .OUT(na1082_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2522_1), .IN6(na1082_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1082_2 ( .OUT(na1082_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1082_1_i) );
// C_MX4b/D///      x93y80     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_1 ( .OUT(na1083_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2520_2), .IN6(na1083_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_2 ( .OUT(na1083_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1083_1_i) );
// C_MX4b/D///      x93y77     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1084_1 ( .OUT(na1084_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1084_1), .IN6(na5593_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1084_2 ( .OUT(na1084_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1084_1_i) );
// C_MX4b/D///      x86y75     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_1 ( .OUT(na1085_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9398_2), .IN6(na5592_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_2 ( .OUT(na1085_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1085_1_i) );
// C_MX4b/D///      x115y111     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1086_1 ( .OUT(na1086_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1086_1), .IN6(na482_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1086_2 ( .OUT(na1086_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1086_1_i) );
// C_MX4b/D///      x119y109     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_1 ( .OUT(na1087_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9236_2),
                      .IN8(na9399_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_2 ( .OUT(na1087_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1087_1_i) );
// C_MX4b/D///      x116y109     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1088_1 ( .OUT(na1088_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na581_1), .IN6(na9401_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1088_2 ( .OUT(na1088_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1088_1_i) );
// C_MX4b/D///      x105y111     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1089_1 ( .OUT(na1089_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1089_1), .IN6(na472_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1089_2 ( .OUT(na1089_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1089_1_i) );
// C_MX4b/D///      x103y109     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1090_1 ( .OUT(na1090_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1090_1), .IN6(na1091_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1090_2 ( .OUT(na1090_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1090_1_i) );
// C_AND////      x93y86     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1091_1 ( .OUT(na1091_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na9404_2), .IN7(na2539_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x107y107     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1092_1 ( .OUT(na1092_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1092_1), .IN6(na961_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1092_2 ( .OUT(na1092_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1092_1_i) );
// C_MX4b/D///      x107y105     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1093_1 ( .OUT(na1093_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1093_1), .IN6(na993_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1093_2 ( .OUT(na1093_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1093_1_i) );
// C_MX4b/D///      x103y107     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1094_1 ( .OUT(na1094_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1095_2),
                      .IN8(na9402_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1094_2 ( .OUT(na1094_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1094_1_i) );
// C_///AND/      x98y77     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1095_4 ( .OUT(na1095_2), .IN1(1'b1), .IN2(~na9404_2), .IN3(na2542_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y105     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1096_1 ( .OUT(na1096_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1096_1),
                      .IN8(na1097_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1096_2 ( .OUT(na1096_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1096_1_i) );
// C_///AND/      x94y78     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1097_4 ( .OUT(na1097_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1113_1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x99y91     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1098_1 ( .OUT(na1098_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1098_1), .IN6(na1099_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1098_2 ( .OUT(na1098_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1098_1_i) );
// C_AND////      x93y88     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1099_1 ( .OUT(na1099_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(~na1113_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x99y111     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1100_1 ( .OUT(na1100_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1100_1), .IN6(na1101_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1100_2 ( .OUT(na1100_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1100_1_i) );
// C_///AND/      x91y82     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1101_4 ( .OUT(na1101_2), .IN1(1'b1), .IN2(na2545_2), .IN3(~na1113_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x105y109     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1102_1 ( .OUT(na1102_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1102_1), .IN6(na1103_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1102_2 ( .OUT(na1102_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1102_1_i) );
// C_AND////      x101y96     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1103_1 ( .OUT(na1103_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(na2547_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x101y109     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1104_1 ( .OUT(na1104_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1104_1), .IN6(na1105_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1104_2 ( .OUT(na1104_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1104_1_i) );
// C_///AND/      x93y90     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1105_4 ( .OUT(na1105_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1113_1), .IN4(na2548_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x103y111     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1106_1 ( .OUT(na1106_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1106_1), .IN6(na991_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1106_2 ( .OUT(na1106_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1106_1_i) );
// C_MX2b////      x129y50     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1108_1 ( .OUT(na1108_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na500_2), .IN5(1'b0), .IN6(~na2972_2), .IN7(1'b0), .IN8(~na7090_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x107y109     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1109_1 ( .OUT(na1109_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1109_1), .IN6(na1110_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1109_2 ( .OUT(na1109_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1109_1_i) );
// C_AND////      x103y96     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1110_1 ( .OUT(na1110_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na9404_2), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x96y95     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_1 ( .OUT(na1111_1_i), .IN1(1'b1), .IN2(na1112_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1111_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_2 ( .OUT(na1111_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1111_1_i) );
// C_///AND/      x97y92     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1112_4 ( .OUT(na1112_2), .IN1(na906_1), .IN2(na1024_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x102y81     80'h00_FE00_80_0000_0C88_2F14
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1113_1 ( .OUT(na1113_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na8_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1113_2 ( .OUT(na1113_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1113_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1113_4 ( .OUT(na1113_2_i), .IN1(~na32_1), .IN2(na467_1), .IN3(~na1113_2), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1113_5 ( .OUT(na1113_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1113_2_i) );
// C_MX4b/D///      x112y99     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1114_1 ( .OUT(na1114_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1114_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1114_2 ( .OUT(na1114_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1114_1_i) );
// C_MX4b/D///      x111y97     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1115_1 ( .OUT(na1115_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1115_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1115_2 ( .OUT(na1115_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1115_1_i) );
// C_MX4b/D///      x110y93     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_1 ( .OUT(na1116_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1116_1),
                      .IN8(na1097_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_2 ( .OUT(na1116_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1116_1_i) );
// C_MX4b/D///      x112y94     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1117_1 ( .OUT(na1117_1_i), .IN1(1'b1), .IN2(~na454_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na1117_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1117_2 ( .OUT(na1117_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1117_1_i) );
// C_MX4b/D///      x114y93     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1118_1 ( .OUT(na1118_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9408_2), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1118_2 ( .OUT(na1118_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1118_1_i) );
// C_MX4b/D///      x122y69     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1119_1 ( .OUT(na1119_1_i), .IN1(na898_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1119_1),
                      .IN8(na1120_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1119_2 ( .OUT(na1119_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1119_1_i) );
// C_AND////      x126y68     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1120_1 ( .OUT(na1120_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3878_2), .IN6(na7044_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x112y98     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_1 ( .OUT(na1121_1_i), .IN1(1'b1), .IN2(~na454_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na1121_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_2 ( .OUT(na1121_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1121_1_i) );
// C_MX4b/D///      x118y97     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1123_1 ( .OUT(na1123_1_i), .IN1(1'b1), .IN2(~na454_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na9410_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1123_2 ( .OUT(na1123_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1123_1_i) );
// C_MX4b/D///      x103y101     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1124_1 ( .OUT(na1124_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1124_1), .IN6(na1099_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1124_2 ( .OUT(na1124_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1124_1_i) );
// C_///AND/D      x69y108     80'h00_F600_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1125_4 ( .OUT(na1125_2_i), .IN1(1'b1), .IN2(na43_2), .IN3(1'b1), .IN4(na404_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1125_5 ( .OUT(na1125_2), .CLK(na4116_1), .EN(~na359_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1125_2_i) );
// C_AND/D//AND/D      x77y99     80'h00_F600_80_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1126_1 ( .OUT(na1126_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3698_1), .IN6(na410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1126_2 ( .OUT(na1126_1), .CLK(na4116_1), .EN(~na56_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1126_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1126_4 ( .OUT(na1126_2_i), .IN1(1'b1), .IN2(na3700_1), .IN3(na9220_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1126_5 ( .OUT(na1126_2), .CLK(na4116_1), .EN(~na56_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1126_2_i) );
// C_AND/D///      x117y79     80'h00_FE00_00_0000_0888_8524
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1127_1 ( .OUT(na1127_1_i), .IN1(~na3256_1), .IN2(na3345_1), .IN3(na4204_2), .IN4(~na6626_1), .IN5(~na3290_1), .IN6(1'b1),
                      .IN7(na3596_2), .IN8(na983_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1127_2 ( .OUT(na1127_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1127_1_i) );
// C_///ORAND/D      x106y86     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1128_4 ( .OUT(na1128_2_i), .IN1(na1129_1), .IN2(na7094_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1128_5 ( .OUT(na1128_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1128_2_i) );
// C_AND////      x109y87     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2922_1), .IN7(na298_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x101y62     80'h00_FE18_00_0000_0888_5CFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1130_1 ( .OUT(na1130_1), .IN1(1'b1), .IN2(na1042_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1131_1), .IN7(~na1132_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1130_5 ( .OUT(na1130_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1130_1) );
// C_AND////      x99y74     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na566_1), .IN6(na435_1), .IN7(na433_2), .IN8(na9230_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y63     80'h00_0018_00_0000_0888_4F15
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1132_1 ( .OUT(na1132_1), .IN1(~na1167_1), .IN2(1'b1), .IN3(~na1165_2), .IN4(~na1134_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na1165_1),
                      .IN8(na1134_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND/D      x110y58     80'h00_FE00_80_0000_0C88_3D3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(na7096_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_2 ( .OUT(na1134_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1134_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1134_4 ( .OUT(na1134_2_i), .IN1(na8130_1), .IN2(~na2998_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1134_5 ( .OUT(na1134_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1134_2_i) );
// C_XOR////      x108y58     80'h00_0018_00_0000_0C66_A300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1130_1), .IN7(na1136_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x102y57     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1136_4 ( .OUT(na1136_2), .IN1(~na2991_1), .IN2(na974_1), .IN3(~na7098_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y53     80'h00_0018_00_0040_0CF6_5300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1), .IN1(1'b1), .IN2(~na4108_2), .IN3(~na3849_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na1130_1), .IN7(~na1136_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x107y87     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1138_1 ( .OUT(na1138_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1139_1), .IN6(na9415_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1138_2 ( .OUT(na1138_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1138_1_i) );
// C_AND////      x97y83     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(~na1113_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x112y88     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7100_1), .IN6(na1141_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_2 ( .OUT(na1140_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1140_1_i) );
// C_AND////      x111y88     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1694_1), .IN6(1'b1), .IN7(na298_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x122y70     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1142_1 ( .OUT(na1142_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7102_2), .IN6(na1143_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1142_2 ( .OUT(na1142_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1142_1_i) );
// C_///AND/      x109y82     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1143_4 ( .OUT(na1143_2), .IN1(1'b1), .IN2(na3125_1), .IN3(na298_1), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x96y105     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_1 ( .OUT(na1145_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1145_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_2 ( .OUT(na1145_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1145_1_i) );
// C_MX4b/D///      x108y108     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9417_2), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_2 ( .OUT(na1147_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1147_1_i) );
// C_MX4b/D///      x112y106     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1148_1 ( .OUT(na1148_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na1148_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1148_2 ( .OUT(na1148_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1148_1_i) );
// C_MX4b/D///      x108y106     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1149_1 ( .OUT(na1149_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na1149_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1149_2 ( .OUT(na1149_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1149_1_i) );
// C_MX4b/D///      x112y104     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1150_1 ( .OUT(na1150_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9419_2), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1150_2 ( .OUT(na1150_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1150_1_i) );
// C_MX4b/D///      x110y108     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_1 ( .OUT(na1151_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na1151_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_2 ( .OUT(na1151_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1151_1_i) );
// C_MX4b/D///      x112y108     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1152_1 ( .OUT(na1152_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na1152_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1152_2 ( .OUT(na1152_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1152_1_i) );
// C_MX4b/D///      x108y105     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1153_1 ( .OUT(na1153_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9421_2), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1153_2 ( .OUT(na1153_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1153_1_i) );
// C_MX4b/D///      x100y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_1 ( .OUT(na1154_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9423_2), .IN6(na1073_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_2 ( .OUT(na1154_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1154_1_i) );
// C_MX4b/D///      x102y94     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_1 ( .OUT(na1155_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na9425_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_2 ( .OUT(na1155_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1155_1_i) );
// C_MX4b/D///      x104y94     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1156_1 ( .OUT(na1156_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9426_2), .IN6(na454_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1156_2 ( .OUT(na1156_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1156_1_i) );
// C_MX4b/D///      x100y94     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_1 ( .OUT(na1157_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9427_2), .IN6(na1078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_2 ( .OUT(na1157_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1157_1_i) );
// C_MX4b/D///      x106y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1158_1 ( .OUT(na1158_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9429_2), .IN6(na893_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1158_2 ( .OUT(na1158_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1158_1_i) );
// C_MX4b/D///      x112y96     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1159_1 ( .OUT(na1159_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9431_2), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1159_2 ( .OUT(na1159_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1159_1_i) );
// C_AND///AND/      x115y100     80'h00_0078_00_0000_0C88_4FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1160_1 ( .OUT(na1160_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1113_1), .IN8(na2530_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1160_4 ( .OUT(na1160_2), .IN1(na428_1), .IN2(1'b1), .IN3(na490_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x116y114     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_1 ( .OUT(na1161_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na833_1),
                      .IN8(na1161_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_2 ( .OUT(na1161_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1161_1_i) );
// C_MX4b/D///      x118y114     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1162_1 ( .OUT(na1162_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9432_2), .IN6(na482_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1162_2 ( .OUT(na1162_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1162_1_i) );
// C_MX4b/D///      x116y112     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_1 ( .OUT(na1163_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9236_2),
                      .IN8(na1163_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_2 ( .OUT(na1163_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1163_1_i) );
// C_MX4b/D///      x116y110     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1164_1 ( .OUT(na1164_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na581_1), .IN6(na9435_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1164_2 ( .OUT(na1164_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1164_1_i) );
// C_ORAND/D//ORAND/D      x110y57     80'h00_FE00_80_0000_0C88_3B3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8132_2), .IN6(~na1166_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_2 ( .OUT(na1165_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1165_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1165_4 ( .OUT(na1165_2_i), .IN1(na8132_1), .IN2(~na3000_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1165_5 ( .OUT(na1165_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1165_2_i) );
// C_MX4a////      x109y52     80'h00_0018_00_0040_0CF9_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1166_1 ( .OUT(na1166_1), .IN1(~na4106_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3847_1), .IN5(1'b1), .IN6(na1130_1), .IN7(~na1136_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x111y59     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1167_1 ( .OUT(na1167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1168_1), .IN6(na7106_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1167_2 ( .OUT(na1167_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1167_1_i) );
// C_ICOMP////      x105y59     80'h00_0018_00_0000_0C88_65FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1167_1), .IN6(1'b0), .IN7(na1136_2), .IN8(~na9411_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x98y62     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1169_1 ( .OUT(na1169_1_i), .IN1(~na9414_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3845_1),
                      .IN8(na1169_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1169_2 ( .OUT(na1169_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1169_1_i) );
// C_MX4b/D///      x98y59     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_1 ( .OUT(na1170_1_i), .IN1(na9414_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1170_1),
                      .IN8(na3843_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_2 ( .OUT(na1170_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1170_1_i) );
// C_MX4b/D///      x99y59     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_1 ( .OUT(na1171_1_i), .IN1(na9414_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9436_2),
                      .IN8(na3843_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_2 ( .OUT(na1171_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1171_1_i) );
// C_MX4b/D///      x94y62     80'h00_FE00_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1172_1 ( .OUT(na1172_1_i), .IN1(na9414_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9437_2),
                      .IN8(~na1172_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1172_2 ( .OUT(na1172_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1172_1_i) );
// C_AND/D///      x85y98     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_1 ( .OUT(na1173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1174_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_2 ( .OUT(na1173_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1173_1_i) );
// C_///AND/      x93y89     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1174_4 ( .OUT(na1174_2), .IN1(na488_1), .IN2(na1131_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND*/D      x94y82     80'h00_FE00_80_0000_0C87_3E77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1175_1 ( .OUT(na1175_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1176_2), .IN6(na7108_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1175_2 ( .OUT(na1175_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1175_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1175_4 ( .OUT(na1175_2_i), .IN1(~na1246_1), .IN2(~na9438_2), .IN3(~na1248_1), .IN4(~na2989_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1175_5 ( .OUT(na1175_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1175_2_i) );
// C_///ORAND/      x87y83     80'h00_0060_00_0000_0C08_FFC7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1176_4 ( .OUT(na1176_2), .IN1(~na1224_1), .IN2(~na1173_1), .IN3(1'b0), .IN4(na1175_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//AND/D      x90y83     80'h00_FE00_80_0000_0C88_3E2F
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1177_1 ( .OUT(na1177_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_2), .IN6(na1179_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1177_2 ( .OUT(na1177_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1177_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1177_4 ( .OUT(na1177_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1177_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1177_5 ( .OUT(na1177_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1177_2_i) );
// C_///ORAND/      x83y85     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1178_4 ( .OUT(na1178_2), .IN1(~na7111_1), .IN2(1'b0), .IN3(~na1177_1), .IN4(na7109_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y82     80'h00_0018_00_0000_0C88_A7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1179_1 ( .OUT(na1179_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1224_1), .IN6(~na1173_1), .IN7(na1177_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x79y92     80'h00_FE18_00_0000_0888_21C8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1181_1 ( .OUT(na1181_1), .IN1(na1126_2), .IN2(na410_1), .IN3(1'b1), .IN4(na1864_2), .IN5(~na1126_1), .IN6(~na1182_1), .IN7(na4853_2),
                      .IN8(~na1864_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1181_5 ( .OUT(na1181_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1181_1) );
// C_AND////      x87y98     80'h00_0018_00_0000_0888_4555
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1182_1 ( .OUT(na1182_1), .IN1(~na1193_2), .IN2(1'b1), .IN3(~na1191_2), .IN4(1'b1), .IN5(~na1193_1), .IN6(1'b1), .IN7(~na1191_1),
                      .IN8(na1188_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x84y90     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1184_1 ( .OUT(na1184_1_i), .IN1(1'b1), .IN2(~na1181_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3854_1),
                      .IN8(na1184_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1184_2 ( .OUT(na1184_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1184_1_i) );
// C_MX4b/D///      x84y87     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1185_1 ( .OUT(na1185_1_i), .IN1(1'b1), .IN2(na1181_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1185_1),
                      .IN8(na3852_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1185_2 ( .OUT(na1185_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1185_1_i) );
// C_MX4b/D///      x86y87     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1186_1 ( .OUT(na1186_1_i), .IN1(1'b1), .IN2(na1181_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1186_1),
                      .IN8(na3852_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1186_2 ( .OUT(na1186_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1186_1_i) );
// C_MX4b/D///      x87y87     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1187_1 ( .OUT(na1187_1_i), .IN1(1'b1), .IN2(na1181_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1187_1), .IN6(~na9442_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1187_2 ( .OUT(na1187_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1187_1_i) );
// C_ORAND/D///      x88y96     80'h00_FE00_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1188_1 ( .OUT(na1188_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7114_2), .IN6(~na1190_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1188_2 ( .OUT(na1188_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1188_1_i) );
// C_///XOR/      x85y94     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1189_4 ( .OUT(na1189_2), .IN1(na1178_2), .IN2(~na1181_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x83y98     80'h00_0018_00_0040_0CF9_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1190_1 ( .OUT(na1190_1), .IN1(~na4113_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na3862_2), .IN5(~na1178_2), .IN6(1'b1), .IN7(na9441_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND/D      x88y95     80'h00_FE00_80_0000_0C88_3B3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1191_1 ( .OUT(na1191_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7122_2), .IN6(~na1192_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1191_2 ( .OUT(na1191_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1191_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1191_4 ( .OUT(na1191_2_i), .IN1(na7122_1), .IN2(na1218_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1191_5 ( .OUT(na1191_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1191_2_i) );
// C_MX4a////      x83y96     80'h00_0018_00_0040_0CF9_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1192_1 ( .OUT(na1192_1), .IN1(~na4113_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3862_1), .IN5(~na1178_2), .IN6(1'b1), .IN7(na9441_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND/D      x89y95     80'h00_FE00_80_0000_0C88_3D3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1193_1 ( .OUT(na1193_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1194_1), .IN6(na7118_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1193_2 ( .OUT(na1193_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1193_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1193_4 ( .OUT(na1193_2_i), .IN1(na7120_2), .IN2(~na1196_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1193_5 ( .OUT(na1193_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1193_2_i) );
// C_MX4a////      x81y95     80'h00_0018_00_0040_0CF6_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1194_1 ( .OUT(na1194_1), .IN1(1'b1), .IN2(~na4111_2), .IN3(~na3860_2), .IN4(1'b1), .IN5(na1178_2), .IN6(1'b1), .IN7(na9441_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x85y96     80'h00_0018_00_0040_0CF6_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1196_1 ( .OUT(na1196_1), .IN1(1'b1), .IN2(~na4111_1), .IN3(~na3860_1), .IN4(1'b1), .IN5(na1178_2), .IN6(1'b1), .IN7(na9441_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x106y112     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1197_1 ( .OUT(na1197_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9443_2), .IN6(na472_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1197_2 ( .OUT(na1197_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1197_1_i) );
// C_MX4b/D///      x106y114     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1198_1 ( .OUT(na1198_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9444_2), .IN6(na1091_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1198_2 ( .OUT(na1198_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1198_1_i) );
// C_MX4b/D///      x110y112     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_1 ( .OUT(na1199_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9446_2), .IN6(na961_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_2 ( .OUT(na1199_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1199_1_i) );
// C_MX4b/D///      x106y108     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1200_1 ( .OUT(na1200_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9448_2), .IN6(na993_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1200_2 ( .OUT(na1200_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1200_1_i) );
// C_MX4b/D///      x106y110     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1201_1 ( .OUT(na1201_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1095_2),
                      .IN8(na1201_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1201_2 ( .OUT(na1201_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1201_1_i) );
// C_MX4b/D///      x102y107     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1202_1 ( .OUT(na1202_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1202_1),
                      .IN8(na1097_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1202_2 ( .OUT(na1202_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1202_1_i) );
// C_MX4b/D///      x104y110     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1203_1 ( .OUT(na1203_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9450_2), .IN6(na1099_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1203_2 ( .OUT(na1203_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1203_1_i) );
// C_MX4b/D///      x100y112     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1204_1 ( .OUT(na1204_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9452_2), .IN6(na1101_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1204_2 ( .OUT(na1204_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1204_1_i) );
// C_MX4b/D///      x102y112     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1205_1 ( .OUT(na1205_1_i), .IN1(~na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1139_1), .IN6(na9453_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1205_2 ( .OUT(na1205_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1205_1_i) );
// C_MX4b/D///      x102y110     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1206_1 ( .OUT(na1206_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9454_2), .IN6(na1103_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1206_2 ( .OUT(na1206_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1206_1_i) );
// C_MX4b/D///      x108y114     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1207_1 ( .OUT(na1207_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9456_2), .IN6(na1105_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1207_2 ( .OUT(na1207_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1207_1_i) );
// C_MX4b/D///      x104y112     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1208_1 ( .OUT(na1208_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9458_2), .IN6(na991_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1208_2 ( .OUT(na1208_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1208_1_i) );
// C_MX4b/D///      x108y112     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1209_1 ( .OUT(na1209_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9459_2), .IN6(na1110_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1209_2 ( .OUT(na1209_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1209_1_i) );
// C_MX4b/D///      x110y110     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1210_1 ( .OUT(na1210_1_i), .IN1(na1034_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9460_2), .IN6(na1211_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1210_2 ( .OUT(na1210_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1210_1_i) );
// C_AND////      x109y100     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1211_1 ( .OUT(na1211_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na9404_2), .IN7(na2551_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x102y76     80'h00_FE00_80_0000_0C08_FF38
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1212_4 ( .OUT(na1212_2_i), .IN1(na906_1), .IN2(na1024_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1212_5 ( .OUT(na1212_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1212_2_i) );
// C_AND/D///      x100y89     80'h00_FE00_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1213_1 ( .OUT(na1213_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1214_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1213_2 ( .OUT(na1213_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1213_1_i) );
// C_MX2a////      x87y86     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1214_1 ( .OUT(na1214_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1213_1), .IN4(~na159_1), .IN5(na9360_2), .IN6(na1024_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x103y93     80'h00_FE00_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1215_1 ( .OUT(na1215_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9361_2), .IN6(na1024_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1215_2 ( .OUT(na1215_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1215_1_i) );
// C_MX4b/D///      x97y113     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1216_1 ( .OUT(na1216_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1216_1), .IN6(na1287_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1216_2 ( .OUT(na1216_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1216_1_i) );
// C_///ICOMP/      x85y92     80'h00_0060_00_0000_0C08_FF56
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1218_4 ( .OUT(na1218_2), .IN1(na1178_2), .IN2(~na1181_1), .IN3(na1191_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x86y80     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1219_1 ( .OUT(na1219_1_i), .IN1(~na1178_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3858_1),
                      .IN8(na1219_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1219_2 ( .OUT(na1219_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1219_1_i) );
// C_MX4b/D///      x88y77     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1220_1 ( .OUT(na1220_1_i), .IN1(na1178_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1220_1),
                      .IN8(na3856_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1220_2 ( .OUT(na1220_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1220_1_i) );
// C_MX4b/D///      x82y71     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1221_1 ( .OUT(na1221_1_i), .IN1(na1178_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1221_1),
                      .IN8(na3856_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1221_2 ( .OUT(na1221_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1221_1_i) );
// C_MX4b/D///      x89y79     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1222_1 ( .OUT(na1222_1_i), .IN1(na1178_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1222_1), .IN6(~na9462_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1222_2 ( .OUT(na1222_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1222_1_i) );
// C_AND/D///      x114y53     80'h00_FE00_00_0000_0C88_C2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1223_1 ( .OUT(na1223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3838_1), .IN6(~na9941_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1223_2 ( .OUT(na1223_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1223_1_i) );
// C_MX4b/D///      x93y95     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1224_1 ( .OUT(na1224_1_i), .IN1(na1174_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1224_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1224_2 ( .OUT(na1224_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1224_1_i) );
// C_MX4b/D///      x91y93     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1225_1 ( .OUT(na1225_1_i), .IN1(na1174_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9464_2),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1225_2 ( .OUT(na1225_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1225_1_i) );
// C_MX4b/D///      x117y114     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1226_1 ( .OUT(na1226_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1291_1), .IN6(na1226_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1226_2 ( .OUT(na1226_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1226_1_i) );
// C_MX4b/D///      x113y116     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1227_1 ( .OUT(na1227_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9465_2),
                      .IN8(na1293_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1227_2 ( .OUT(na1227_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1227_1_i) );
// C_MX4b/D///      x117y112     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1228_1 ( .OUT(na1228_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1295_1),
                      .IN8(na9466_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1228_2 ( .OUT(na1228_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1228_1_i) );
// C_MX4b/D///      x115y114     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1229_1 ( .OUT(na1229_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9467_2), .IN6(na1297_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1229_2 ( .OUT(na1229_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1229_1_i) );
// C_MX4b/D///      x121y114     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1230_1 ( .OUT(na1230_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1299_1), .IN6(na1230_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1230_2 ( .OUT(na1230_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1230_1_i) );
// C_MX4b/D///      x119y118     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1231_1 ( .OUT(na1231_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1301_1), .IN6(na1231_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1231_2 ( .OUT(na1231_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1231_1_i) );
// C_MX4b/D///      x109y92     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1232_1 ( .OUT(na1232_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1303_1),
                      .IN8(na9468_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1232_2 ( .OUT(na1232_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1232_1_i) );
// C_MX4b/D///      x119y122     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1233_1 ( .OUT(na1233_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9469_2), .IN6(na2664_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1233_2 ( .OUT(na1233_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1233_1_i) );
// C_MX4b/D///      x121y120     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1234_1 ( .OUT(na1234_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2662_1),
                      .IN8(na9470_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1234_2 ( .OUT(na1234_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1234_1_i) );
// C_MX2a////      x91y90     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1236_1 ( .OUT(na1236_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2681_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1237_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y94     80'h00_0018_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1237_1 ( .OUT(na1237_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9231_2), .IN6(na435_1), .IN7(na436_1), .IN8(~na452_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x115y120     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1238_1 ( .OUT(na1238_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9471_2),
                      .IN8(na1308_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1238_2 ( .OUT(na1238_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1238_1_i) );
// C_MX4b/D///      x117y118     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_1 ( .OUT(na1239_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1310_1), .IN6(na1239_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_2 ( .OUT(na1239_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1239_1_i) );
// C_MX4b/D///      x121y118     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1240_1 ( .OUT(na1240_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1316_1), .IN6(na1240_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1240_2 ( .OUT(na1240_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1240_1_i) );
// C_MX4b/D///      x119y120     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1241_1 ( .OUT(na1241_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9472_2), .IN6(na2659_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1241_2 ( .OUT(na1241_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1241_1_i) );
// C_MX4b/D///      x117y120     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1242_1 ( .OUT(na1242_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1318_1),
                      .IN8(na9473_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1242_2 ( .OUT(na1242_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1242_1_i) );
// C_MX4b/D///      x119y114     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1243_1 ( .OUT(na1243_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9474_2),
                      .IN8(na1323_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1243_2 ( .OUT(na1243_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1243_1_i) );
// C_MX4b/D///      x117y116     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1244_1 ( .OUT(na1244_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1325_1), .IN6(na1244_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1244_2 ( .OUT(na1244_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1244_1_i) );
// C_MX4b/D///      x111y114     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1245_1 ( .OUT(na1245_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9475_2), .IN6(na1327_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1245_2 ( .OUT(na1245_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1245_1_i) );
// C_MX4b/D///      x97y95     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1246_1 ( .OUT(na1246_1_i), .IN1(na1247_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1246_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1246_2 ( .OUT(na1246_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1246_1_i) );
// C_///AND/      x97y81     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1247_4 ( .OUT(na1247_2), .IN1(1'b1), .IN2(na1131_1), .IN3(na567_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x94y89     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1248_1 ( .OUT(na1248_1_i), .IN1(na1247_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1248_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1248_2 ( .OUT(na1248_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1248_1_i) );
// C_AND/D///      x125y52     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1249_1 ( .OUT(na1249_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3796_1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1249_2 ( .OUT(na1249_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1249_1_i) );
// C_AND/D//AND/D      x125y50     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1250_1 ( .OUT(na1250_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3793_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1250_2 ( .OUT(na1250_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1250_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1250_4 ( .OUT(na1250_2_i), .IN1(na3793_1), .IN2(1'b1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1250_5 ( .OUT(na1250_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1250_2_i) );
// C_AND/D//AND/D      x123y49     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1252_1 ( .OUT(na1252_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3791_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1252_2 ( .OUT(na1252_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1252_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1252_4 ( .OUT(na1252_2_i), .IN1(1'b1), .IN2(na3791_1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1252_5 ( .OUT(na1252_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1252_2_i) );
// C_AND/D//AND*/D      x124y48     80'h00_FE00_80_0000_0C87_CAC5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1254_1 ( .OUT(na1254_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3789_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1254_2 ( .OUT(na1254_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1254_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1254_4 ( .OUT(na1254_2_i), .IN1(~na3789_1), .IN2(1'b1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1254_5 ( .OUT(na1254_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1254_2_i) );
// C_AND*/D//AND*/D      x123y47     80'h00_FE00_80_0000_0387_C3C3
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1256_1 ( .OUT(na1256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3787_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1256_2 ( .OUT(na1256_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1256_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1256_4 ( .OUT(na1256_2_i), .IN1(1'b1), .IN2(~na3787_1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1256_5 ( .OUT(na1256_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1256_2_i) );
// C_AND/D//AND*/D      x123y50     80'h00_FE00_80_0000_0C87_CAC5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1258_1 ( .OUT(na1258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3785_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1258_2 ( .OUT(na1258_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1258_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1258_4 ( .OUT(na1258_2_i), .IN1(~na3785_1), .IN2(1'b1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1258_5 ( .OUT(na1258_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1258_2_i) );
// C_AND/D//AND*/D      x124y46     80'h00_FE00_80_0000_0C87_CCC3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1260_1 ( .OUT(na1260_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3782_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1260_2 ( .OUT(na1260_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1260_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1260_4 ( .OUT(na1260_2_i), .IN1(1'b1), .IN2(~na3782_1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1260_5 ( .OUT(na1260_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1260_2_i) );
// C_MX4b/D///      x107y118     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1261_1 ( .OUT(na1261_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9477_2),
                      .IN8(na2244_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1261_2 ( .OUT(na1261_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1261_1_i) );
// C_MX4b/D///      x111y116     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1262_1 ( .OUT(na1262_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2242_1),
                      .IN8(na9478_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1262_2 ( .OUT(na1262_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1262_1_i) );
// C_MX4b/D///      x95y92     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1263_1 ( .OUT(na1263_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9479_2), .IN6(na1329_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1263_2 ( .OUT(na1263_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1263_1_i) );
// C_MX4b/D///      x99y94     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1264_1 ( .OUT(na1264_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2240_1), .IN6(na1264_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1264_2 ( .OUT(na1264_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1264_1_i) );
// C_MX4b/D///      x106y96     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1265_1 ( .OUT(na1265_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2237_1),
                      .IN8(na1265_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1265_2 ( .OUT(na1265_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1265_1_i) );
// C_MX4b/D///      x107y98     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1266_1 ( .OUT(na1266_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9481_2),
                      .IN8(na1331_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1266_2 ( .OUT(na1266_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1266_1_i) );
// C_MX4b/D///      x109y94     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1267_1 ( .OUT(na1267_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2235_1),
                      .IN8(na9482_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1267_2 ( .OUT(na1267_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1267_1_i) );
// C_MX4b/D///      x111y100     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1268_1 ( .OUT(na1268_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9483_2),
                      .IN8(na2166_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1268_2 ( .OUT(na1268_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1268_1_i) );
// C_MX4b/D///      x105y116     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1269_1 ( .OUT(na1269_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9484_2), .IN6(na2161_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1269_2 ( .OUT(na1269_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1269_1_i) );
// C_MX4b/D///      x105y114     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1270_1 ( .OUT(na1270_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2159_1), .IN6(na1270_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1270_2 ( .OUT(na1270_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1270_1_i) );
// C_MX4b/D///      x103y116     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_1 ( .OUT(na1271_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1335_1), .IN6(na1271_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_2 ( .OUT(na1271_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1271_1_i) );
// C_MX4b/D///      x111y118     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1272_1 ( .OUT(na1272_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1340_1),
                      .IN8(na9485_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1272_2 ( .OUT(na1272_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1272_1_i) );
// C_MX4b/D///      x115y118     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1273_1 ( .OUT(na1273_1_i), .IN1(~na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1901_1), .IN6(na1273_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1273_2 ( .OUT(na1273_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1273_1_i) );
// C_ORAND/D///      x99y89     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1274_1 ( .OUT(na1274_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1286_2), .IN6(na7124_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1274_2 ( .OUT(na1274_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1274_1_i) );
// C_AND////      x108y99     80'h00_0018_00_0000_0888_1484
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1275_1 ( .OUT(na1275_1), .IN1(~na1335_1), .IN2(na1284_1), .IN3(na1279_1), .IN4(na1285_1), .IN5(~na1901_1), .IN6(na1284_2),
                      .IN7(~na1340_1), .IN8(~na1289_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y95     80'h00_0018_00_0000_0888_5184
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1279_1 ( .OUT(na1279_1), .IN1(~na1299_1), .IN2(na1282_1), .IN3(na1283_2), .IN4(na1281_2), .IN5(~na1301_1), .IN6(~na1297_1),
                      .IN7(~na1303_1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y96     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1281_4 ( .OUT(na1281_2), .IN1(~na1291_1), .IN2(~na1287_1), .IN3(~na1295_1), .IN4(~na1293_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y96     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1282_1 ( .OUT(na1282_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1316_1), .IN6(~na2659_1), .IN7(~na1318_1),
                      .IN8(~na1323_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y97     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1283_4 ( .OUT(na1283_2), .IN1(~na1310_1), .IN2(~na2664_1), .IN3(~na2662_1), .IN4(~na1308_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y98     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1284_1 ( .OUT(na1284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2240_1), .IN6(~na1329_1), .IN7(~na2237_1),
                      .IN8(~na1331_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1284_4 ( .OUT(na1284_2), .IN1(~na2159_1), .IN2(~na2161_1), .IN3(~na2235_1), .IN4(~na2166_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y96     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1285_1 ( .OUT(na1285_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1325_1), .IN6(~na1327_1), .IN7(~na2242_1),
                      .IN8(~na2244_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x101y89     80'h00_0060_00_0000_0C08_FF7A
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1286_4 ( .OUT(na1286_2), .IN1(na1274_1), .IN2(1'b0), .IN3(~na1111_1), .IN4(~na1212_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x97y100     80'h00_FE00_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1287_1 ( .OUT(na1287_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1030_1),
                      .IN8(~na1288_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1287_2 ( .OUT(na1287_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1287_1_i) );
// C_MX2a////      x104y100     80'h00_0018_00_0040_0C8A_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1288_1 ( .OUT(na1288_1), .IN1(1'b0), .IN2(na1287_1), .IN3(1'b0), .IN4(~na9416_2), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y98     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_1 ( .OUT(na1289_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1032_1), .IN6(~na1290_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_2 ( .OUT(na1289_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1289_1_i) );
// C_MX2a////      x103y94     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1290_1 ( .OUT(na1290_1), .IN1(1'b0), .IN2(~na3999_1), .IN3(1'b0), .IN4(~na1147_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y97     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1291_1 ( .OUT(na1291_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1035_1), .IN6(~na1292_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1291_2 ( .OUT(na1291_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1291_1_i) );
// C_MX2a////      x103y90     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1292_1 ( .OUT(na1292_1), .IN1(1'b0), .IN2(~na3999_2), .IN3(1'b0), .IN4(~na1148_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x102y98     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1293_1 ( .OUT(na1293_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2670_1), .IN6(~na1294_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1293_2 ( .OUT(na1293_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1293_1_i) );
// C_MX2a////      x103y100     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1294_1 ( .OUT(na1294_1), .IN1(~na4013_1), .IN2(1'b0), .IN3(~na9418_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x102y97     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1295_1 ( .OUT(na1295_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1068_1), .IN6(~na1296_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1295_2 ( .OUT(na1295_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1295_1_i) );
// C_MX2a////      x103y102     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1296_1 ( .OUT(na1296_1), .IN1(~na4013_2), .IN2(1'b0), .IN3(~na9420_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y98     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1297_1 ( .OUT(na1297_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1069_1), .IN6(~na1298_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1297_2 ( .OUT(na1297_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1297_1_i) );
// C_MX2a////      x107y102     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1298_1 ( .OUT(na1298_1), .IN1(1'b0), .IN2(~na4015_1), .IN3(1'b0), .IN4(~na1151_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x99y95     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1299_1 ( .OUT(na1299_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1070_1), .IN6(~na1300_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1299_2 ( .OUT(na1299_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1299_1_i) );
// C_MX2a////      x93y104     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1300_1 ( .OUT(na1300_1), .IN1(1'b0), .IN2(~na4015_2), .IN3(1'b0), .IN4(~na1152_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y99     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1301_1 ( .OUT(na1301_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1071_1), .IN6(~na1302_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1301_2 ( .OUT(na1301_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1301_1_i) );
// C_MX2a////      x113y108     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1302_1 ( .OUT(na1302_1), .IN1(~na4017_1), .IN2(1'b0), .IN3(~na1153_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y99     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1303_1 ( .OUT(na1303_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1072_1), .IN6(~na1304_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1303_2 ( .OUT(na1303_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1303_1_i) );
// C_MX2a////      x107y104     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1304_1 ( .OUT(na1304_1), .IN1(~na4017_2), .IN2(1'b0), .IN3(~na1154_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x91y87     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1306_1 ( .OUT(na1306_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1314_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1307_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y86     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1307_4 ( .OUT(na1307_2), .IN1(na9229_2), .IN2(na435_1), .IN3(na433_2), .IN4(~na452_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x102y100     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_1 ( .OUT(na1308_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1077_1), .IN6(~na1309_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_2 ( .OUT(na1308_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1308_1_i) );
// C_MX2a////      x107y100     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1309_1 ( .OUT(na1309_1), .IN1(~na3990_1), .IN2(1'b0), .IN3(~na9428_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x111y99     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1310_1 ( .OUT(na1310_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1080_1), .IN6(~na1311_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1310_2 ( .OUT(na1310_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1310_1_i) );
// C_MX2a////      x103y110     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1311_1 ( .OUT(na1311_1), .IN1(~na3990_2), .IN2(1'b0), .IN3(~na1158_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x96y93     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1312_1 ( .OUT(na1312_1_i), .IN1(1'b1), .IN2(na1313_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1312_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1312_2 ( .OUT(na1312_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1312_1_i) );
// C_AND////      x97y86     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na906_1), .IN6(na459_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x90y97     80'h00_FE00_80_0000_0C88_3335
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1314_1 ( .OUT(na1314_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1315_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1314_2 ( .OUT(na1314_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1314_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1314_4 ( .OUT(na1314_2_i), .IN1(~na1306_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1314_5 ( .OUT(na1314_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1314_2_i) );
// C_MX2a////      x115y76     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1315_1 ( .OUT(na1315_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1314_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1307_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y101     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1316_1 ( .OUT(na1316_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2669_1), .IN6(~na1317_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1316_2 ( .OUT(na1316_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1316_1_i) );
// C_MX2a////      x105y102     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1317_1 ( .OUT(na1317_1), .IN1(1'b0), .IN2(~na3992_1), .IN3(1'b0), .IN4(~na1159_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x112y101     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1318_1 ( .OUT(na1318_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1086_1), .IN6(~na1319_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1318_2 ( .OUT(na1318_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1318_1_i) );
// C_MX2a////      x103y106     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1319_1 ( .OUT(na1319_1), .IN1(~na3994_1), .IN2(1'b0), .IN3(~na9433_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y85     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1321_1 ( .OUT(na1321_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2677_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1322_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y82     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1322_1 ( .OUT(na1322_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9229_2), .IN6(na435_1), .IN7(na433_1), .IN8(~na452_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x118y120     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_1 ( .OUT(na1323_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1087_1), .IN6(~na1324_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_2 ( .OUT(na1323_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1323_1_i) );
// C_MX2a////      x113y106     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1324_1 ( .OUT(na1324_1), .IN1(~na3994_2), .IN2(1'b0), .IN3(~na9434_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x115y119     80'h00_FE00_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_1 ( .OUT(na1325_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1088_1),
                      .IN8(~na1326_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_2 ( .OUT(na1325_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1325_1_i) );
// C_MX2a////      x108y104     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1326_1 ( .OUT(na1326_1), .IN1(1'b0), .IN2(~na3996_1), .IN3(1'b0), .IN4(~na1164_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x105y118     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1327_1 ( .OUT(na1327_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1089_1), .IN6(~na1328_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1327_2 ( .OUT(na1327_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1327_1_i) );
// C_MX2a////      x107y106     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1328_1 ( .OUT(na1328_1), .IN1(1'b0), .IN2(~na3996_2), .IN3(1'b0), .IN4(~na1197_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x101y102     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1329_1 ( .OUT(na1329_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1093_1), .IN6(~na1330_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1329_2 ( .OUT(na1329_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1329_1_i) );
// C_MX2a////      x109y104     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1330_1 ( .OUT(na1330_1), .IN1(1'b0), .IN2(~na4001_1), .IN3(1'b0), .IN4(~na1200_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x102y102     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1331_1 ( .OUT(na1331_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1098_1), .IN6(~na1332_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1331_2 ( .OUT(na1331_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1331_1_i) );
// C_MX2a////      x105y108     80'h00_0018_00_0040_0C55_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1332_1 ( .OUT(na1332_1), .IN1(~na4003_2), .IN2(1'b0), .IN3(~na9451_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x122y72     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1_i), .IN1(~na898_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1334_1),
                      .IN8(na1333_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1333_2 ( .OUT(na1333_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1333_1_i) );
// C_AND////      x126y65     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1334_1 ( .OUT(na1334_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3878_1), .IN6(na7044_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x99y103     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1335_1 ( .OUT(na1335_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1106_1), .IN6(~na1336_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1335_2 ( .OUT(na1335_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1335_1_i) );
// C_MX2a////      x105y104     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1336_1 ( .OUT(na1336_1), .IN1(1'b0), .IN2(~na4009_1), .IN3(1'b0), .IN4(~na1208_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x90y95     80'h00_FE00_80_0000_0C88_1F35
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1337_1 ( .OUT(na1337_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1338_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1337_2 ( .OUT(na1337_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1337_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1337_4 ( .OUT(na1337_2_i), .IN1(~na1877_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1337_5 ( .OUT(na1337_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1337_2_i) );
// C_MX2a////      x92y91     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1338_1 ( .OUT(na1338_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1337_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1339_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y84     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1339_1 ( .OUT(na1339_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9226_2), .IN6(na435_2), .IN7(na436_1), .IN8(~na452_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y103     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1340_1 ( .OUT(na1340_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1109_1), .IN6(~na1341_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1340_2 ( .OUT(na1340_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1340_1_i) );
// C_MX2a////      x111y104     80'h00_0018_00_0040_0CAA_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1341_1 ( .OUT(na1341_1), .IN1(1'b0), .IN2(~na4009_2), .IN3(1'b0), .IN4(~na1209_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x117y101     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1342_1 ( .OUT(na1342_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1342_1), .IN6(na482_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1342_2 ( .OUT(na1342_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1342_1_i) );
// C_AND/D//AND/D      x51y110     80'h00_FE00_80_0000_0C88_AAF2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1343_1 ( .OUT(na1343_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3816_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1343_2 ( .OUT(na1343_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1343_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1343_4 ( .OUT(na1343_2_i), .IN1(na971_1), .IN2(~na1343_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1343_5 ( .OUT(na1343_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1343_2_i) );
// C_///AND/D      x96y89     80'h00_FE00_80_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1344_4 ( .OUT(na1344_2_i), .IN1(~na1345_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1344_5 ( .OUT(na1344_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1344_2_i) );
// C_MX2a////      x87y99     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1344_2), .IN4(~na159_1), .IN5(na853_2), .IN6(na564_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x90y98     80'h00_FE00_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1346_1 ( .OUT(na1346_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1347_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1346_2 ( .OUT(na1346_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1346_1_i) );
// C_MX2a////      x89y97     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1347_1 ( .OUT(na1347_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na9491_2), .IN4(~na159_1), .IN5(na906_1), .IN6(na564_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x100y88     80'h00_FE00_80_0000_0C08_FF38
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1349_4 ( .OUT(na1349_2_i), .IN1(na853_2), .IN2(na564_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1349_5 ( .OUT(na1349_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1349_2_i) );
// C_MX4b/D///      x95y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1350_1 ( .OUT(na1350_1_i), .IN1(na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1350_1), .IN6(na5179_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1350_2 ( .OUT(na1350_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1350_1_i) );
// C_AND/D///      x97y92     80'h00_FE00_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_1 ( .OUT(na1351_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1352_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_2 ( .OUT(na1351_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1351_1_i) );
// C_MX2a////      x96y87     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1352_1 ( .OUT(na1352_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na9492_2), .IN4(~na159_1), .IN5(na9266_2), .IN6(na564_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x98y94     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_1 ( .OUT(na1353_1_i), .IN1(na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9493_2), .IN6(na5179_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_2 ( .OUT(na1353_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1353_1_i) );
// C_MX4b/D///      x91y111     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1354_1 ( .OUT(na1354_1_i), .IN1(na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1354_1), .IN6(na5181_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1354_2 ( .OUT(na1354_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1354_1_i) );
// C_AND/D//AND/D      x74y73     80'h00_FE00_80_0000_0C88_3335
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1355_1 ( .OUT(na1355_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1356_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1355_2 ( .OUT(na1355_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1355_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1355_4 ( .OUT(na1355_2_i), .IN1(~na2684_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1355_5 ( .OUT(na1355_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1355_2_i) );
// C_MX2a////      x87y78     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1356_1 ( .OUT(na1356_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1355_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1357_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y74     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1357_4 ( .OUT(na1357_2), .IN1(na566_1), .IN2(na435_2), .IN3(na436_1), .IN4(~na9228_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x69y102     80'h00_FE00_00_0000_0C88_2AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1358_1 ( .OUT(na1358_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na4069_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1358_2 ( .OUT(na1358_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1358_1_i) );
// C_AND/D//AND/D      x74y75     80'h00_FE00_80_0000_0C88_1F1F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_1 ( .OUT(na1359_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1360_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_2 ( .OUT(na1359_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1359_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1359_4 ( .OUT(na1359_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na2686_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1359_5 ( .OUT(na1359_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1359_2_i) );
// C_MX2a////      x90y89     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1360_1 ( .OUT(na1360_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1359_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1361_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y84     80'h00_0018_00_0000_0C88_82FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1361_1 ( .OUT(na1361_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na566_1), .IN6(~na435_1), .IN7(na433_1), .IN8(na9230_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x91y109     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1362_1 ( .OUT(na1362_1_i), .IN1(na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1362_1), .IN6(na5183_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1362_2 ( .OUT(na1362_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1362_1_i) );
// C_MX4b/D///      x89y109     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_1 ( .OUT(na1363_1_i), .IN1(na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1363_1), .IN6(na5183_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_2 ( .OUT(na1363_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1363_1_i) );
// C_MX4b/D///      x96y106     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1_i), .IN1(~na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na1364_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_2 ( .OUT(na1364_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1364_1_i) );
// C_AND*/D//AND*/D      x124y45     80'h00_FE00_80_0000_0387_C5C5
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1365_1 ( .OUT(na1365_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3780_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1365_2 ( .OUT(na1365_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1365_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1365_4 ( .OUT(na1365_2_i), .IN1(~na3780_1), .IN2(1'b1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1365_5 ( .OUT(na1365_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1365_2_i) );
// C_MX4b/D///      x96y104     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_1 ( .OUT(na1366_1_i), .IN1(~na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na1366_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_2 ( .OUT(na1366_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1366_1_i) );
// C_MX4b/D///      x116y82     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1367_1 ( .OUT(na1367_1_i), .IN1(1'b1), .IN2(~na981_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9862_2),
                      .IN8(na1367_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1367_2 ( .OUT(na1367_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1367_1_i) );
// C_AND///AND/      x65y89     80'h00_0078_00_0000_0C88_C4F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1370_1 ( .OUT(na1370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na714_1), .IN6(na1462_2), .IN7(1'b1), .IN8(na503_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1370_4 ( .OUT(na1370_2), .IN1(na714_2), .IN2(~na504_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x111y84     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1371_1 ( .OUT(na1371_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9499_2), .IN6(na3050_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1371_2 ( .OUT(na1371_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1371_1_i) );
// C_AND/D///      x65y79     80'h00_FE00_00_0000_0888_2F2C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1372_1 ( .OUT(na1372_1_i), .IN1(1'b1), .IN2(na397_2), .IN3(na403_1), .IN4(~na406_1), .IN5(1'b1), .IN6(1'b1), .IN7(na517_2),
                      .IN8(~na42_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1372_2 ( .OUT(na1372_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1372_1_i) );
// C_///AND/D      x77y79     80'h00_FE00_80_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1373_4 ( .OUT(na1373_2_i), .IN1(1'b1), .IN2(na2172_2), .IN3(na542_1), .IN4(na3319_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1373_5 ( .OUT(na1373_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1373_2_i) );
// C_AND/D//AND*/D      x123y44     80'h00_FE00_80_0000_0C87_CAC5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1375_1 ( .OUT(na1375_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3776_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1375_2 ( .OUT(na1375_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1375_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1375_4 ( .OUT(na1375_2_i), .IN1(~na3776_1), .IN2(1'b1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1375_5 ( .OUT(na1375_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1375_2_i) );
// C_AND/D///      x58y78     80'h00_FE00_00_0000_0C88_2AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1377_1 ( .OUT(na1377_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na514_2), .IN6(1'b1), .IN7(na403_1), .IN8(~na1378_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1377_2 ( .OUT(na1377_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1377_1_i) );
// C_MX2b////      x54y80     80'h00_0018_00_0040_0AA8_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1378_1 ( .OUT(na1378_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na347_2), .IN4(1'b1), .IN5(1'b0), .IN6(na9202_2), .IN7(1'b0), .IN8(~na1377_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x66y93     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1379_4 ( .OUT(na1379_2_i), .IN1(1'b1), .IN2(na7129_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1379_5 ( .OUT(na1379_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1379_2_i) );
// C_AND////      x70y86     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1380_1 ( .OUT(na1380_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9815_2), .IN6(na504_1), .IN7(na359_1), .IN8(na3324_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y94     80'h00_0018_00_0040_0A55_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1381_1 ( .OUT(na1381_1), .IN1(na9324_2), .IN2(1'b1), .IN3(na359_2), .IN4(1'b1), .IN5(~na1388_1), .IN6(1'b0), .IN7(~na1379_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x112y90     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1382_1 ( .OUT(na1382_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9501_2), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1382_2 ( .OUT(na1382_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1382_1_i) );
// C_ORAND/D///      x65y74     80'h00_FA00_00_0000_0C88_73FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1383_1 ( .OUT(na1383_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na7131_1), .IN7(~na1384_1),
                      .IN8(~na1385_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1383_2 ( .OUT(na1383_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1383_1_i) );
// C_MX2a////      x80y69     80'h00_0018_00_0040_0CCC_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1384_1 ( .OUT(na1384_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2558_1), .IN4(~na9206_2), .IN5(~na2555_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x72y70     80'h00_0060_00_0000_0C0E_FF3C
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1385_4 ( .OUT(na1385_2), .IN1(1'b0), .IN2(na7132_2), .IN3(1'b0), .IN4(~na2556_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x74y71     80'h00_FE00_80_0000_0C88_A8FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1372_1), .IN6(na9215_2), .IN7(na1387_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1387_2 ( .OUT(na1387_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1387_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1387_4 ( .OUT(na1387_2_i), .IN1(1'b1), .IN2(na5985_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1387_5 ( .OUT(na1387_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1387_2_i) );
// C_AND/D///      x65y83     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1388_1 ( .OUT(na1388_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na7134_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1388_2 ( .OUT(na1388_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1388_1_i) );
// C_MX2a////      x53y125     80'h00_0018_00_0040_0C55_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1389_1 ( .OUT(na1389_1), .IN1(~na7135_1), .IN2(1'b0), .IN3(~na1379_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na731_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x123y74     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1390_4 ( .OUT(na1390_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7136_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1390_5 ( .OUT(na1390_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1390_2_i) );
// C_AND/D///      x75y105     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1392_1 ( .OUT(na1392_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1), .IN8(na7140_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1392_2 ( .OUT(na1392_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1392_1_i) );
// C_MX4a////D      x59y108     80'h00_FA18_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1393_1 ( .OUT(na1393_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b0), .IN4(~na1395_1), .IN5(1'b1), .IN6(na5953_2), .IN7(~na2316_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1393_5 ( .OUT(na1393_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1393_1) );
// C_AND////      x68y114     80'h00_0018_00_0000_0888_5238
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1395_1 ( .OUT(na1395_1), .IN1(na7141_2), .IN2(na7145_1), .IN3(1'b1), .IN4(~na7146_2), .IN5(na7141_1), .IN6(~na7142_2), .IN7(~na7144_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x72y90     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1399_4 ( .OUT(na1399_2_i), .IN1(1'b1), .IN2(na7147_1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1399_5 ( .OUT(na1399_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1399_2_i) );
// C_AND////      x70y85     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1400_1 ( .OUT(na1400_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9245_2), .IN6(na3317_1), .IN7(na359_1), .IN8(na3324_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x122y73     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1401_4 ( .OUT(na1401_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7148_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1401_5 ( .OUT(na1401_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1401_2_i) );
// C_ORAND*/D///      x61y91     80'h00_FE00_00_0000_0788_AFE3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1403_1 ( .OUT(na1403_1_i), .IN1(1'b0), .IN2(~na7152_1), .IN3(na7154_1), .IN4(na731_1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1403_2 ( .OUT(na1403_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1403_1_i) );
// C_ORAND*/D///      x53y123     80'h00_FE00_00_0000_0788_AFE3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1405_1 ( .OUT(na1405_1_i), .IN1(1'b0), .IN2(~na7152_1), .IN3(na7157_2), .IN4(na731_1), .IN5(1'b1), .IN6(1'b1), .IN7(na403_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1405_2 ( .OUT(na1405_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1405_1_i) );
// C_AND/D///      x68y90     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1407_1 ( .OUT(na1407_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9216_2), .IN6(1'b1), .IN7(na7158_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1407_2 ( .OUT(na1407_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1407_1_i) );
// C_AND/D///      x76y89     80'h00_FE00_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1408_1 ( .OUT(na1408_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9201_2), .IN6(na716_1), .IN7(na403_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1408_2 ( .OUT(na1408_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1408_1_i) );
// C_ORAND*/D///      x120y63     80'h00_FE00_00_0000_0788_BF3E
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1409_1 ( .OUT(na1409_1_i), .IN1(na2991_1), .IN2(na9365_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na7160_1),
                      .IN8(~na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1409_2 ( .OUT(na1409_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1409_1_i) );
// C_MX4b/D///      x113y90     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_1 ( .OUT(na1411_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9504_2),
                      .IN8(na3052_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_2 ( .OUT(na1411_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1411_1_i) );
// C_///AND/D      x117y71     80'h00_FE00_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1412_4 ( .OUT(na1412_2_i), .IN1(1'b1), .IN2(~na7161_1), .IN3(1'b1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1412_5 ( .OUT(na1412_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1412_2_i) );
// C_///AND/D      x75y112     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1414_4 ( .OUT(na1414_2_i), .IN1(na9216_2), .IN2(1'b1), .IN3(na6381_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1414_5 ( .OUT(na1414_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1414_2_i) );
// C_AND/D///      x110y78     80'h00_FE00_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1415_1 ( .OUT(na1415_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(~na7165_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1415_2 ( .OUT(na1415_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1415_1_i) );
// C_///AND/      x97y87     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1416_4 ( .OUT(na1416_2), .IN1(na7078_1), .IN2(na435_1), .IN3(na9265_2), .IN4(~na452_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x112y77     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1418_1 ( .OUT(na1418_1_i), .IN1(na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1418_1),
                      .IN8(na6478_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1418_2 ( .OUT(na1418_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1418_1_i) );
// C_AND/D///      x107y70     80'h00_F900_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1419_1 ( .OUT(na1419_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6118_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2829_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1419_2 ( .OUT(na1419_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1419_1_i) );
// C_///AND/D      x103y81     80'h00_FE00_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1420_4 ( .OUT(na1420_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1421_1), .IN4(~na7171_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1420_5 ( .OUT(na1420_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1420_2_i) );
// C_AND////      x102y69     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1421_1 ( .OUT(na1421_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9954_2), .IN6(~na435_1), .IN7(na433_2), .IN8(~na1055_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y50     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1425_4 ( .OUT(na1425_2), .IN1(na6118_2), .IN2(1'b1), .IN3(na7176_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x119y41     80'h00_F900_80_0000_0C88_CCC5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1427_1 ( .OUT(na1427_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4064_1), .IN7(1'b1), .IN8(na1425_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1427_2 ( .OUT(na1427_1), .CLK(~na4116_1), .EN(na3254_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1427_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1427_4 ( .OUT(na1427_2_i), .IN1(~na1427_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1425_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1427_5 ( .OUT(na1427_2), .CLK(~na4116_1), .EN(na3254_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1427_2_i) );
// C_AND/D//AND/D      x120y40     80'h00_F900_80_0000_0C88_CACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1429_1 ( .OUT(na1429_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4066_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1425_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1429_2 ( .OUT(na1429_1), .CLK(~na4116_1), .EN(na3254_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1429_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1429_4 ( .OUT(na1429_2_i), .IN1(1'b1), .IN2(na4064_2), .IN3(1'b1), .IN4(na1425_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1429_5 ( .OUT(na1429_2), .CLK(~na4116_1), .EN(na3254_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1429_2_i) );
// C_AND/D///      x117y41     80'h00_F900_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1430_1 ( .OUT(na1430_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4066_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1425_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1430_2 ( .OUT(na1430_1), .CLK(~na4116_1), .EN(na3254_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1430_1_i) );
// C_///AND/D      x115y71     80'h00_FE00_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1431_4 ( .OUT(na1431_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1421_1), .IN4(~na7178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1431_5 ( .OUT(na1431_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1431_2_i) );
// C_AND/D//AND/D      x76y113     80'h00_FE00_80_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1433_1 ( .OUT(na1433_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9216_2), .IN6(1'b1), .IN7(na6381_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1433_2 ( .OUT(na1433_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1433_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1433_4 ( .OUT(na1433_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na6380_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1433_5 ( .OUT(na1433_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1433_2_i) );
// C_///AND/      x89y99     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1434_4 ( .OUT(na1434_2), .IN1(~na9809_2), .IN2(~na3299_2), .IN3(~na3301_1), .IN4(~na3216_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x106y88     80'h00_FE00_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1435_1 ( .OUT(na1435_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1436_1), .IN6(1'b0), .IN7(na7183_1), .IN8(~na7182_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1435_2 ( .OUT(na1435_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1435_1_i) );
// C_AND////      x103y83     80'h00_0018_00_0000_0C88_32FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1436_1 ( .OUT(na1436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(~na435_1), .IN7(1'b1), .IN8(~na452_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x102y90     80'h00_FE00_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1438_1 ( .OUT(na1438_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1436_1), .IN6(1'b0), .IN7(na7185_1), .IN8(~na7184_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1438_2 ( .OUT(na1438_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1438_1_i) );
// C_ORAND/D///      x112y85     80'h00_FE00_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1441_1 ( .OUT(na1441_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1436_1), .IN6(1'b0), .IN7(na7187_1), .IN8(~na7186_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1441_2 ( .OUT(na1441_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1441_1_i) );
// C_///ORAND/D      x104y85     80'h00_FE00_80_0000_0C08_FFBA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1443_4 ( .OUT(na1443_2_i), .IN1(na1436_1), .IN2(1'b0), .IN3(na7189_1), .IN4(~na7188_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1443_5 ( .OUT(na1443_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1443_2_i) );
// C_MX4b/D///      x114y86     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1445_1 ( .OUT(na1445_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na457_1), .IN6(~na1446_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1445_2 ( .OUT(na1445_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1445_1_i) );
// C_MX2b////      x115y88     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1446_1 ( .OUT(na1446_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9302_2), .IN8(~na4037_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y86     80'h00_0018_00_0000_0888_4184
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1447_1 ( .OUT(na1447_1), .IN1(~na3034_1), .IN2(na1451_1), .IN3(na1457_2), .IN4(na1456_1), .IN5(~na3040_1), .IN6(~na3038_1),
                      .IN7(~na3036_1), .IN8(na1456_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y86     80'h00_0018_00_0000_0888_1238
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1), .IN1(na1455_1), .IN2(na1453_1), .IN3(1'b1), .IN4(~na3052_1), .IN5(na1454_2), .IN6(~na3050_1), .IN7(~na3056_1),
                      .IN8(~na3054_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y88     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1453_1 ( .OUT(na1453_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3044_1), .IN6(~na3046_1), .IN7(~na3042_1),
                      .IN8(~na3048_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y85     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1454_4 ( .OUT(na1454_2), .IN1(~na3081_1), .IN2(~na3077_1), .IN3(~na3068_1), .IN4(~na3079_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y85     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1455_1 ( .OUT(na1455_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3058_1), .IN6(~na3060_1), .IN7(~na3062_1),
                      .IN8(~na1445_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x114y84     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1456_1 ( .OUT(na1456_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3093_1), .IN6(~na3091_1), .IN7(~na3097_1),
                      .IN8(~na3095_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1456_4 ( .OUT(na1456_2), .IN1(~na3099_1), .IN2(~na3105_1), .IN3(~na3103_1), .IN4(~na3101_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y85     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1457_4 ( .OUT(na1457_2), .IN1(~na3089_1), .IN2(~na3085_1), .IN3(~na3083_1), .IN4(~na3087_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x111y87     80'h00_FE00_00_0000_0C88_DAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1458_1 ( .OUT(na1458_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1436_1), .IN6(1'b0), .IN7(~na7190_1), .IN8(na7191_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1458_2 ( .OUT(na1458_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1458_1_i) );
// C_///AND/D      x106y76     80'h00_FE00_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1460_4 ( .OUT(na1460_2_i), .IN1(na1436_1), .IN2(1'b1), .IN3(~na7192_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1460_5 ( .OUT(na1460_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1460_2_i) );
// C_ORAND/D//ORAND/D      x65y90     80'h00_FE00_80_0000_0C88_AEAE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1462_1 ( .OUT(na1462_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1370_2), .IN6(na1463_2), .IN7(na403_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1462_2 ( .OUT(na1462_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1462_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1462_4 ( .OUT(na1462_2_i), .IN1(na1370_1), .IN2(na713_1), .IN3(na403_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1462_5 ( .OUT(na1462_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1462_2_i) );
// C_///AND/      x71y82     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1463_4 ( .OUT(na1463_2), .IN1(~na9201_2), .IN2(na716_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x106y82     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1464_4 ( .OUT(na1464_2_i), .IN1(na1436_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na7198_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1464_5 ( .OUT(na1464_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1464_2_i) );
// C_AND////      x116y108     80'h00_0018_00_0000_0888_54F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1467_1 ( .OUT(na1467_1), .IN1(~na7202_2), .IN2(na7203_2), .IN3(1'b1), .IN4(1'b1), .IN5(~na7204_1), .IN6(na7203_1), .IN7(~na7206_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x100y79     80'h00_FE00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1470_4 ( .OUT(na1470_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1471_1), .IN4(na2695_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1470_5 ( .OUT(na1470_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1470_2_i) );
// C_AND////      x102y79     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1471_1 ( .OUT(na1471_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9954_2), .IN6(na435_2), .IN7(~na9227_2),
                      .IN8(na9223_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x101y75     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1473_4 ( .OUT(na1473_2_i), .IN1(na2697_1), .IN2(1'b1), .IN3(na1471_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1473_5 ( .OUT(na1473_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1473_2_i) );
// C_AND/D///      x94y88     80'h00_FE00_00_0000_0888_3358
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1475_1 ( .OUT(na1475_1_i), .IN1(na9954_2), .IN2(na435_2), .IN3(~na9227_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na7208_1), .IN7(1'b1),
                      .IN8(~na1476_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1475_2 ( .OUT(na1475_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1475_1_i) );
// C_MX2b////      x100y74     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1476_1 ( .OUT(na1476_1), .IN1(1'b1), .IN2(~na1042_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na9660_2), .IN6(~na6592_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x91y86     80'h00_FE00_00_0000_0888_AAB3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1479_1 ( .OUT(na1479_1_i), .IN1(1'b0), .IN2(~na435_1), .IN3(na7210_1), .IN4(~na7209_1), .IN5(na9954_2), .IN6(1'b0), .IN7(na433_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1479_2 ( .OUT(na1479_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1479_1_i) );
// C_AND/D//AND/D      x74y104     80'h00_FE00_80_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1481_1 ( .OUT(na1481_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7211_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1481_2 ( .OUT(na1481_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1481_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1481_4 ( .OUT(na1481_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na7133_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1481_5 ( .OUT(na1481_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1481_2_i) );
// C_AND/D///      x114y71     80'h00_FE00_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1482_1 ( .OUT(na1482_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1421_1), .IN8(~na7212_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1482_2 ( .OUT(na1482_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1482_1_i) );
// C_///AND/D      x113y71     80'h00_FE00_80_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1484_4 ( .OUT(na1484_2_i), .IN1(1'b1), .IN2(~na7216_1), .IN3(na1421_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1484_5 ( .OUT(na1484_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1484_2_i) );
// C_AND/D///      x109y71     80'h00_FE00_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1486_1 ( .OUT(na1486_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1421_1), .IN8(~na7220_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1486_2 ( .OUT(na1486_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1486_1_i) );
// C_///AND/D      x110y70     80'h00_FE00_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1488_4 ( .OUT(na1488_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1421_1), .IN4(~na7224_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1488_5 ( .OUT(na1488_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1488_2_i) );
// C_AND/D///      x116y77     80'h00_FE00_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1490_1 ( .OUT(na1490_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na7228_1), .IN7(na1421_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1490_2 ( .OUT(na1490_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1490_1_i) );
// C_AND/D///      x72y83     80'h00_FE00_00_0000_0C88_83FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1492_1 ( .OUT(na1492_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1493_1), .IN7(na403_1), .IN8(na503_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1492_2 ( .OUT(na1492_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1492_1_i) );
// C_MX2b////      x81y80     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1493_1 ( .OUT(na1493_1), .IN1(1'b1), .IN2(~na343_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1492_1), .IN8(~na9209_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x74y100     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1494_1 ( .OUT(na1494_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3925_2), .IN8(~na1495_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1494_5 ( .OUT(na1494_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1494_1) );
// C_MX2b////      x62y106     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1495_1 ( .OUT(na1495_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3958_1), .IN8(na1496_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y114     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1496_1 ( .OUT(na1496_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2225_1), .IN7(1'b0), .IN8(~na689_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x68y95     80'h00_FE00_80_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1497_1 ( .OUT(na1497_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7232_1), .IN6(1'b1), .IN7(na403_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1497_2 ( .OUT(na1497_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1497_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1497_4 ( .OUT(na1497_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na403_1), .IN4(na7025_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1497_5 ( .OUT(na1497_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1497_2_i) );
// C_MX2b////D      x80y95     80'h00_F618_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1498_1 ( .OUT(na1498_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1499_1), .IN8(na3923_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1498_5 ( .OUT(na1498_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1498_1) );
// C_MX2b////      x72y109     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1499_1 ( .OUT(na1499_1), .IN1(1'b1), .IN2(na397_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1500_1), .IN6(~na5848_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x59y113     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1500_1 ( .OUT(na1500_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na731_1), .IN5(1'b0), .IN6(~na2219_1), .IN7(1'b0), .IN8(~na674_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x78y91     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1502_1 ( .OUT(na1502_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3916_1), .IN8(~na1503_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1502_5 ( .OUT(na1502_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1502_1) );
// C_MX2b////      x72y104     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1503_1 ( .OUT(na1503_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na5842_1), .IN8(na1504_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x60y110     80'h00_0018_00_0040_0CAA_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1504_1 ( .OUT(na1504_1), .IN1(1'b0), .IN2(~na2207_1), .IN3(1'b0), .IN4(~na629_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na731_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x108y71     80'h00_FE00_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1506_4 ( .OUT(na1506_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1421_1), .IN4(~na7235_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1506_5 ( .OUT(na1506_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1506_2_i) );
// C_AND/D///      x105y72     80'h00_FE00_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1509_1 ( .OUT(na1509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7240_1), .IN6(1'b1), .IN7(na1421_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1509_2 ( .OUT(na1509_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1509_1_i) );
// C_MX4b/D///      x120y96     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1512_1 ( .OUT(na1512_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9516_2), .IN6(na893_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1512_2 ( .OUT(na1512_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1512_1_i) );
// C_AND////      x89y70     80'h00_0018_00_0000_0888_3448
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1524_1 ( .OUT(na1524_1), .IN1(na1045_2), .IN2(na1525_2), .IN3(~na66_1), .IN4(na61_1), .IN5(~na86_1), .IN6(na1525_1), .IN7(1'b1),
                      .IN8(~na37_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y76     80'h00_0078_00_0000_0C88_AC45
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1525_1 ( .OUT(na1525_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1525_2), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1525_4 ( .OUT(na1525_2), .IN1(~na32_1), .IN2(1'b1), .IN3(~na1113_1), .IN4(na9134_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y76     80'h00_0018_00_0000_0888_3825
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1527_1 ( .OUT(na1527_1), .IN1(~na86_1), .IN2(1'b1), .IN3(na66_1), .IN4(~na61_1), .IN5(na1045_2), .IN6(na1525_2), .IN7(1'b1),
                      .IN8(~na1046_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x92y75     80'h00_0018_00_0000_0888_CB3A
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1530_1 ( .OUT(na1530_1), .IN1(na1045_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na37_1), .IN5(na6828_1), .IN6(~na1525_2), .IN7(1'b0),
                      .IN8(na9518_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y74     80'h00_0018_00_0000_0888_3845
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1531_1 ( .OUT(na1531_1), .IN1(~na86_1), .IN2(1'b1), .IN3(~na66_1), .IN4(na61_1), .IN5(na1045_2), .IN6(na1525_2), .IN7(1'b1),
                      .IN8(~na1046_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x110y70     80'h00_FE00_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1532_1 ( .OUT(na1532_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na7266_1), .IN7(na1421_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1532_2 ( .OUT(na1532_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1532_1_i) );
// C_AND/D///      x110y68     80'h00_FE00_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1535_1 ( .OUT(na1535_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1421_1), .IN8(~na7271_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1535_2 ( .OUT(na1535_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1535_1_i) );
// C_///AND/D      x102y75     80'h00_FE00_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1538_4 ( .OUT(na1538_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1421_1), .IN4(~na7276_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1538_5 ( .OUT(na1538_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1538_2_i) );
// C_AND/D///      x97y90     80'h00_FE00_00_0000_0C88_21FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1542_1 ( .OUT(na1542_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7282_1), .IN6(~na435_1), .IN7(na7210_2),
                      .IN8(~na452_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1542_2 ( .OUT(na1542_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1542_1_i) );
// C_///AND/D      x95y88     80'h00_FE00_80_0000_0C08_FF14
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1545_4 ( .OUT(na1545_2_i), .IN1(~na9226_2), .IN2(na435_2), .IN3(~na7286_1), .IN4(~na452_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1545_5 ( .OUT(na1545_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1545_2_i) );
// C_///ORAND/D      x118y69     80'h00_FE00_80_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1548_4 ( .OUT(na1548_2_i), .IN1(1'b0), .IN2(na874_1), .IN3(~na7290_1), .IN4(na7291_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1548_5 ( .OUT(na1548_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1548_2_i) );
// C_///ORAND/D      x106y73     80'h00_FE00_80_0000_0C08_FFBC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1550_4 ( .OUT(na1550_2_i), .IN1(1'b0), .IN2(na874_1), .IN3(na7293_1), .IN4(~na7292_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1550_5 ( .OUT(na1550_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1550_2_i) );
// C_MX2b////D      x75y81     80'h00_F618_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1552_1 ( .OUT(na1552_1), .IN1(1'b1), .IN2(~na727_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3933_2), .IN8(~na1553_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1552_5 ( .OUT(na1552_2), .CLK(na4116_1), .EN(~na711_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1552_1) );
// C_MX2b////      x66y102     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1553_1 ( .OUT(na1553_1), .IN1(1'b1), .IN2(~na397_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3968_1), .IN8(na1554_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y112     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1554_1 ( .OUT(na1554_1), .IN1(1'b1), .IN2(~na9325_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2185_1), .IN6(~na582_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x67y94     80'h00_FE00_80_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1555_1 ( .OUT(na1555_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7294_1), .IN7(na403_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1555_2 ( .OUT(na1555_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1555_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1555_4 ( .OUT(na1555_2_i), .IN1(na6999_1), .IN2(1'b1), .IN3(na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1555_5 ( .OUT(na1555_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1555_2_i) );
// C_///ORAND/D      x111y67     80'h00_FE00_80_0000_0C08_FFBC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1556_4 ( .OUT(na1556_2_i), .IN1(1'b0), .IN2(na874_1), .IN3(na7296_1), .IN4(~na7295_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1556_5 ( .OUT(na1556_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1556_2_i) );
// C_///ORAND/D      x116y66     80'h00_FE00_80_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1558_4 ( .OUT(na1558_2_i), .IN1(1'b0), .IN2(na874_1), .IN3(~na7297_2), .IN4(na7298_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1558_5 ( .OUT(na1558_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1558_2_i) );
// C_///ORAND/D      x112y66     80'h00_FE00_80_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1560_4 ( .OUT(na1560_2_i), .IN1(1'b0), .IN2(na874_1), .IN3(~na7299_2), .IN4(na7300_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1560_5 ( .OUT(na1560_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1560_2_i) );
// C_///AND/D      x119y61     80'h00_FE00_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1562_4 ( .OUT(na1562_2_i), .IN1(1'b1), .IN2(na874_1), .IN3(1'b1), .IN4(~na7301_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1562_5 ( .OUT(na1562_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1562_2_i) );
// C_///AND/D      x118y63     80'h00_FE00_80_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1564_4 ( .OUT(na1564_2_i), .IN1(~na7305_1), .IN2(na874_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1564_5 ( .OUT(na1564_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1564_2_i) );
// C_///AND/D      x95y90     80'h00_FE00_80_0000_0C08_FF21
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1568_4 ( .OUT(na1568_2_i), .IN1(~na9232_2), .IN2(~na435_1), .IN3(na433_1), .IN4(~na7313_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1568_5 ( .OUT(na1568_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1568_2_i) );
// C_///ORAND/D      x98y92     80'h00_FE00_80_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1571_4 ( .OUT(na1571_2_i), .IN1(1'b0), .IN2(na565_2), .IN3(~na7317_1), .IN4(na7318_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1571_5 ( .OUT(na1571_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1571_2_i) );
// C_ORAND/D///      x98y89     80'h00_FE00_00_0000_0C88_BCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1573_1 ( .OUT(na1573_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na565_2), .IN7(na7320_2), .IN8(~na7319_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1573_2 ( .OUT(na1573_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1573_1_i) );
// C_ORAND/D///      x98y90     80'h00_FE00_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1575_1 ( .OUT(na1575_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na565_2), .IN7(~na7321_1), .IN8(na7322_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1575_2 ( .OUT(na1575_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1575_1_i) );
// C_///ORAND/D      x97y83     80'h00_FE00_80_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1577_4 ( .OUT(na1577_2_i), .IN1(1'b0), .IN2(na565_2), .IN3(~na7323_1), .IN4(na7324_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1577_5 ( .OUT(na1577_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1577_2_i) );
// C_///ORAND/D      x100y86     80'h00_FE00_80_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1579_4 ( .OUT(na1579_2_i), .IN1(1'b0), .IN2(na565_2), .IN3(~na7325_1), .IN4(na7326_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1579_5 ( .OUT(na1579_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1579_2_i) );
// C_MX4a////D      x58y104     80'h00_FA18_00_0040_0CB3_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1583_1 ( .OUT(na1583_1), .IN1(~na1584_1), .IN2(~na5953_1), .IN3(1'b0), .IN4(1'b1), .IN5(na1586_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na9912_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1583_5 ( .OUT(na1583_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1583_1) );
// C_ORAND////      x63y113     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1584_1 ( .OUT(na1584_1), .IN1(~na3313_2), .IN2(~na2211_1), .IN3(~na5476_2), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                      .IN8(~na1587_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y73     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1586_1 ( .OUT(na1586_1), .IN1(na3264_1), .IN2(1'b1), .IN3(~na3265_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9900_2),
                      .IN8(na5961_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x58y92     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1587_1 ( .OUT(na1587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7334_1), .IN7(na403_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1587_2 ( .OUT(na1587_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1587_1_i) );
// C_///AND/D      x86y96     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1590_4 ( .OUT(na1590_2_i), .IN1(na7339_1), .IN2(na565_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1590_5 ( .OUT(na1590_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1590_2_i) );
// C_///AND/      x91y78     80'h00_0060_00_0000_0C08_FF12
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1595_4 ( .OUT(na1595_2), .IN1(na1045_2), .IN2(~na64_1), .IN3(~na9160_2), .IN4(~na1046_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x89y75     80'h00_FE00_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1597_1 ( .OUT(na1597_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(na1598_1), .IN7(1'b1), .IN8(na9117_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1597_2 ( .OUT(na1597_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1597_1_i) );
// C_AND////      x91y76     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1598_1 ( .OUT(na1598_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na566_1), .IN6(na435_1), .IN7(na433_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x97y74     80'h00_FE00_80_0000_0C88_C82F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_1 ( .OUT(na1599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(na1598_1), .IN7(1'b1), .IN8(na9118_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_2 ( .OUT(na1599_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1599_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1599_4 ( .OUT(na1599_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1421_1), .IN4(~na7245_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1599_5 ( .OUT(na1599_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1599_2_i) );
// C_MX4a////D      x52y102     80'h00_FA18_00_0040_0CB3_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1600_1 ( .OUT(na1600_1), .IN1(~na1601_1), .IN2(~na5953_1), .IN3(1'b0), .IN4(1'b1), .IN5(na1603_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na9912_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1600_5 ( .OUT(na1600_2), .CLK(na4116_1), .EN(na3244_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1600_1) );
// C_ORAND////      x59y109     80'h00_0018_00_0000_0888_7F77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1601_1 ( .OUT(na1601_1), .IN1(~na3313_2), .IN2(~na2205_1), .IN3(~na5473_1), .IN4(~na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3308_1),
                      .IN8(~na1604_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y63     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1603_1 ( .OUT(na1603_1), .IN1(~na3264_1), .IN2(1'b1), .IN3(na3265_1), .IN4(1'b1), .IN5(na5958_1), .IN6(na5280_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x62y122     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1604_1 ( .OUT(na1604_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9216_2), .IN6(1'b1), .IN7(na7353_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1604_2 ( .OUT(na1604_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1604_1_i) );
// C_AND/D//AND/D      x98y73     80'h00_FE00_80_0000_0C88_A82F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1605_1 ( .OUT(na1605_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(na1598_1), .IN7(na9119_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1605_2 ( .OUT(na1605_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1605_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1605_4 ( .OUT(na1605_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1421_1), .IN4(~na7250_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1605_5 ( .OUT(na1605_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1605_2_i) );
// C_AND/D//AND/D      x96y73     80'h00_FE00_80_0000_0C88_A8A3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1606_1 ( .OUT(na1606_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(na1598_1), .IN7(na9120_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1606_2 ( .OUT(na1606_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1606_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1606_4 ( .OUT(na1606_2_i), .IN1(1'b1), .IN2(~na7255_1), .IN3(na1421_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1606_5 ( .OUT(na1606_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1606_2_i) );
// C_AND/D//AND/D      x95y73     80'h00_FE00_80_0000_0C88_C8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1607_1 ( .OUT(na1607_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(na1598_1), .IN7(1'b1), .IN8(na9121_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1607_2 ( .OUT(na1607_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1607_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1607_4 ( .OUT(na1607_2_i), .IN1(1'b1), .IN2(na7260_1), .IN3(na1421_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1607_5 ( .OUT(na1607_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1607_2_i) );
// C_AND////      x85y70     80'h00_0018_00_0000_0888_3428
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1612_1 ( .OUT(na1612_1), .IN1(na1045_2), .IN2(na1525_2), .IN3(na66_1), .IN4(~na61_1), .IN5(~na86_1), .IN6(na1525_1), .IN7(1'b1),
                      .IN8(~na37_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y70     80'h00_0018_00_0000_0C88_18FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1614_1 ( .OUT(na1614_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1045_2), .IN6(na69_1), .IN7(~na9160_2), .IN8(~na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x105y80     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1616_1 ( .OUT(na1616_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7363_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1616_2 ( .OUT(na1616_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1616_1_i) );
// C_///AND/D      x100y78     80'h00_FE00_80_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1618_4 ( .OUT(na1618_2_i), .IN1(na1416_2), .IN2(~na7367_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1618_5 ( .OUT(na1618_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1618_2_i) );
// C_AND/D///      x59y89     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1620_1 ( .OUT(na1620_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7371_1), .IN7(na403_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1620_2 ( .OUT(na1620_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1620_1_i) );
// C_///AND/D      x103y84     80'h00_FE00_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1621_4 ( .OUT(na1621_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(~na7372_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1621_5 ( .OUT(na1621_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1621_2_i) );
// C_MX4b/D///      x104y78     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1623_1 ( .OUT(na1623_1_i), .IN1(na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9527_2), .IN6(na6477_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1623_2 ( .OUT(na1623_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1623_1_i) );
// C_AND/D///      x106y81     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1624_1 ( .OUT(na1624_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7376_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1624_2 ( .OUT(na1624_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1624_1_i) );
// C_///ORAND*/D      x67y82     80'h00_F600_80_0000_0C07_FFC7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1626_4 ( .OUT(na1626_2_i), .IN1(~na5930_1), .IN2(~na43_1), .IN3(1'b0), .IN4(na42_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1626_5 ( .OUT(na1626_2), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1626_2_i) );
// C_AND/D///      x103y89     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1627_1 ( .OUT(na1627_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7381_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1627_2 ( .OUT(na1627_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1627_1_i) );
// C_///AND/D      x105y92     80'h00_FE00_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1629_4 ( .OUT(na1629_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(~na7385_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1629_5 ( .OUT(na1629_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1629_2_i) );
// C_AND/D///      x103y81     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1631_1 ( .OUT(na1631_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1631_2 ( .OUT(na1631_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1631_1_i) );
// C_///AND/D      x106y78     80'h00_FE00_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1633_4 ( .OUT(na1633_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(~na7393_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1633_5 ( .OUT(na1633_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1633_2_i) );
// C_///AND/D      x108y83     80'h00_FE00_80_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1635_4 ( .OUT(na1635_2_i), .IN1(na1416_2), .IN2(~na7397_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1635_5 ( .OUT(na1635_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1635_2_i) );
// C_AND/D///      x109y82     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1637_1 ( .OUT(na1637_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7401_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1637_2 ( .OUT(na1637_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1637_1_i) );
// C_AND/D///      x100y78     80'h00_FE00_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1639_1 ( .OUT(na1639_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(~na7405_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1639_2 ( .OUT(na1639_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1639_1_i) );
// C_///AND/D      x109y83     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1641_4 ( .OUT(na1641_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na7409_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1641_5 ( .OUT(na1641_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1641_2_i) );
// C_AND/D///      x107y80     80'h00_FE00_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1643_1 ( .OUT(na1643_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(~na7413_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1643_2 ( .OUT(na1643_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1643_1_i) );
// C_///AND/D      x106y83     80'h00_FE00_80_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1645_4 ( .OUT(na1645_2_i), .IN1(na1416_2), .IN2(~na7417_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1645_5 ( .OUT(na1645_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1645_2_i) );
// C_///AND/D      x107y79     80'h00_FE00_80_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1647_4 ( .OUT(na1647_2_i), .IN1(~na7421_1), .IN2(1'b1), .IN3(na9505_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1647_5 ( .OUT(na1647_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1647_2_i) );
// C_///AND/D      x105y90     80'h00_FE00_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1649_4 ( .OUT(na1649_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(~na7425_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1649_5 ( .OUT(na1649_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1649_2_i) );
// C_AND/D///      x113y82     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1651_1 ( .OUT(na1651_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7429_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1651_2 ( .OUT(na1651_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1651_1_i) );
// C_MX4b/D///      x125y63     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1653_1 ( .OUT(na1653_1_i), .IN1(na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1653_1), .IN6(na6479_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1653_2 ( .OUT(na1653_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1653_1_i) );
// C_AND/D///      x110y82     80'h00_FE00_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1654_1 ( .OUT(na1654_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(~na7433_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1654_2 ( .OUT(na1654_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1654_1_i) );
// C_MX4b/D///      x97y102     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1656_1 ( .OUT(na1656_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3742_2),
                      .IN8(na9528_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1656_2 ( .OUT(na1656_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1656_1_i) );
// C_MX4b/D///      x119y75     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1658_1 ( .OUT(na1658_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na9529_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1658_2 ( .OUT(na1658_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1658_1_i) );
// C_AND/D///      x108y82     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1659_1 ( .OUT(na1659_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7437_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1659_2 ( .OUT(na1659_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1659_1_i) );
// C_///AND/D      x108y79     80'h00_FE00_80_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1661_4 ( .OUT(na1661_2_i), .IN1(na1416_2), .IN2(~na7441_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1661_5 ( .OUT(na1661_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1661_2_i) );
// C_AND/D///      x108y79     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1663_1 ( .OUT(na1663_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7445_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1663_2 ( .OUT(na1663_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1663_1_i) );
// C_///AND/D      x104y84     80'h00_FE00_80_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1665_4 ( .OUT(na1665_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(~na7449_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1665_5 ( .OUT(na1665_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1665_2_i) );
// C_AND/D///      x107y89     80'h00_FE00_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1667_1 ( .OUT(na1667_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(~na7453_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1667_2 ( .OUT(na1667_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1667_1_i) );
// C_///AND/D      x112y81     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1669_4 ( .OUT(na1669_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na7457_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1669_5 ( .OUT(na1669_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1669_2_i) );
// C_///AND/D      x109y75     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1677_4 ( .OUT(na1677_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na7473_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1677_5 ( .OUT(na1677_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1677_2_i) );
// C_AND/D//AND/D      x103y78     80'h00_FE00_80_0000_0C88_5A3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1679_1 ( .OUT(na1679_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(~na7477_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1679_2 ( .OUT(na1679_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1679_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1679_4 ( .OUT(na1679_2_i), .IN1(1'b1), .IN2(na565_2), .IN3(1'b1), .IN4(~na7327_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1679_5 ( .OUT(na1679_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1679_2_i) );
// C_AND/D//AND/D      x108y77     80'h00_FE00_80_0000_0C88_3A5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1681_1 ( .OUT(na1681_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na7481_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1681_2 ( .OUT(na1681_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1681_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1681_4 ( .OUT(na1681_2_i), .IN1(1'b1), .IN2(na565_2), .IN3(~na7335_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1681_5 ( .OUT(na1681_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1681_2_i) );
// C_AND/D//AND/D      x107y74     80'h00_FE00_80_0000_0C88_F28F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1683_1 ( .OUT(na1683_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1416_2), .IN6(~na1684_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1683_2 ( .OUT(na1683_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1683_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1683_4 ( .OUT(na1683_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na945_1), .IN4(na947_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1683_5 ( .OUT(na1683_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1683_2_i) );
// C_AND////      x95y80     80'h00_0018_00_0000_0888_8811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1684_1 ( .OUT(na1684_1), .IN1(~na7486_2), .IN2(~na7490_2), .IN3(~na7488_2), .IN4(~na7492_2), .IN5(na7487_2), .IN6(na7489_1),
                      .IN7(na7485_1), .IN8(na7491_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x116y75     80'h00_FE00_80_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1689_4 ( .OUT(na1689_2_i), .IN1(~na7493_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1689_5 ( .OUT(na1689_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1689_2_i) );
// C_AND/D///      x108y71     80'h00_FE00_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1691_1 ( .OUT(na1691_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7497_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1691_2 ( .OUT(na1691_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1691_1_i) );
// C_MX4b/D///      x123y80     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1693_1 ( .OUT(na1693_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9530_2),
                      .IN8(na3054_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1693_2 ( .OUT(na1693_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1693_1_i) );
// C_MX4b/D///      x123y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1694_1 ( .OUT(na1694_1_i), .IN1(na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1694_1), .IN6(na6483_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1694_2 ( .OUT(na1694_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1694_1_i) );
// C_MX4b/D///      x93y101     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1695_1 ( .OUT(na1695_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9531_2),
                      .IN8(na3748_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1695_2 ( .OUT(na1695_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1695_1_i) );
// C_MX4b/D///      x119y77     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1697_1 ( .OUT(na1697_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1697_1), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1697_2 ( .OUT(na1697_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1697_1_i) );
// C_///AND/D      x117y72     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1698_4 ( .OUT(na1698_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7501_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1698_5 ( .OUT(na1698_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1698_2_i) );
// C_AND/D///      x117y73     80'h00_FE00_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1700_1 ( .OUT(na1700_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7505_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1700_2 ( .OUT(na1700_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1700_1_i) );
// C_///AND/D      x115y74     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1702_4 ( .OUT(na1702_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7509_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1702_5 ( .OUT(na1702_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1702_2_i) );
// C_///AND/D      x114y73     80'h00_FE00_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1704_4 ( .OUT(na1704_2_i), .IN1(1'b1), .IN2(na9384_2), .IN3(1'b1), .IN4(~na7513_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1704_5 ( .OUT(na1704_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1704_2_i) );
// C_///AND/D      x115y72     80'h00_FE00_80_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1706_4 ( .OUT(na1706_2_i), .IN1(~na7517_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1706_5 ( .OUT(na1706_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1706_2_i) );
// C_AND/D///      x99y75     80'h00_FE00_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1708_1 ( .OUT(na1708_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na7521_1), .IN7(1'b1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1708_2 ( .OUT(na1708_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1708_1_i) );
// C_///AND/D      x115y73     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1710_4 ( .OUT(na1710_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7525_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1710_5 ( .OUT(na1710_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1710_2_i) );
// C_AND/D///      x113y75     80'h00_FE00_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1712_1 ( .OUT(na1712_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7529_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1712_2 ( .OUT(na1712_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1712_1_i) );
// C_///AND/D      x117y75     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1714_4 ( .OUT(na1714_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7533_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1714_5 ( .OUT(na1714_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1714_2_i) );
// C_///AND/D      x117y74     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1716_4 ( .OUT(na1716_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7537_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1716_5 ( .OUT(na1716_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1716_2_i) );
// C_///AND/D      x112y72     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1718_4 ( .OUT(na1718_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7541_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1718_5 ( .OUT(na1718_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1718_2_i) );
// C_AND/D///      x118y74     80'h00_FE00_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1720_1 ( .OUT(na1720_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7545_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1720_2 ( .OUT(na1720_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1720_1_i) );
// C_///AND/D      x126y74     80'h00_FE00_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1722_4 ( .OUT(na1722_2_i), .IN1(1'b1), .IN2(~na7549_1), .IN3(1'b1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1722_5 ( .OUT(na1722_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1722_2_i) );
// C_AND/D///      x117y75     80'h00_FE00_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1724_1 ( .OUT(na1724_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7553_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1724_2 ( .OUT(na1724_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1724_1_i) );
// C_MX4b/D///      x123y89     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1726_1 ( .OUT(na1726_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na581_1), .IN6(na9532_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1726_2 ( .OUT(na1726_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1726_1_i) );
// C_MX4b/D///      x118y64     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1727_1 ( .OUT(na1727_1_i), .IN1(~na1728_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1729_2),
                      .IN8(na1727_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1727_2 ( .OUT(na1727_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1727_1_i) );
// C_AND////      x117y65     80'h00_0018_00_0000_0888_A443
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1728_1 ( .OUT(na1728_1), .IN1(1'b1), .IN2(~na3356_1), .IN3(~na9798_2), .IN4(na841_2), .IN5(~na3594_1), .IN6(na3343_1), .IN7(na3219_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x122y57     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1729_4 ( .OUT(na1729_2), .IN1(~na1730_1), .IN2(1'b1), .IN3(na3885_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x117y63     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1730_1 ( .OUT(na1730_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3180_1), .IN6(1'b1), .IN7(na2163_1), .IN8(na1727_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x125y74     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1731_4 ( .OUT(na1731_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7557_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1731_5 ( .OUT(na1731_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1731_2_i) );
// C_///AND/D      x119y73     80'h00_FE00_80_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1733_4 ( .OUT(na1733_2_i), .IN1(~na7561_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1733_5 ( .OUT(na1733_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1733_2_i) );
// C_AND/D///      x117y74     80'h00_FE00_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1735_1 ( .OUT(na1735_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na7565_1), .IN7(1'b1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1735_2 ( .OUT(na1735_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1735_1_i) );
// C_AND/D///      x115y74     80'h00_FE00_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1737_1 ( .OUT(na1737_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7569_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1737_2 ( .OUT(na1737_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1737_1_i) );
// C_///AND/D      x119y74     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1739_4 ( .OUT(na1739_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na7573_1), .IN4(na1054_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1739_5 ( .OUT(na1739_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1739_2_i) );
// C_AND/D///      x113y71     80'h00_FE00_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1741_1 ( .OUT(na1741_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na9383_2), .IN8(~na7577_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1741_2 ( .OUT(na1741_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1741_1_i) );
// C_AND/D//AND/D      x113y78     80'h00_FE00_80_0000_0C88_4F5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1743_1 ( .OUT(na1743_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7581_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1743_2 ( .OUT(na1743_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1743_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1743_4 ( .OUT(na1743_2_i), .IN1(na1416_2), .IN2(1'b1), .IN3(~na7461_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1743_5 ( .OUT(na1743_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1743_2_i) );
// C_AND/D//AND/D      x111y79     80'h00_FE00_80_0000_0C88_4FF2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1745_1 ( .OUT(na1745_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7585_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1745_2 ( .OUT(na1745_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1745_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1745_4 ( .OUT(na1745_2_i), .IN1(na1416_2), .IN2(~na7465_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1745_5 ( .OUT(na1745_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1745_2_i) );
// C_AND/D//AND/D      x113y74     80'h00_FE00_80_0000_0C88_4FF2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1747_1 ( .OUT(na1747_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7589_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1747_2 ( .OUT(na1747_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1747_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1747_4 ( .OUT(na1747_2_i), .IN1(na1416_2), .IN2(~na7469_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1747_5 ( .OUT(na1747_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1747_2_i) );
// C_AND/D//AND/D      x99y85     80'h00_FE00_80_0000_0C88_4F3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1749_1 ( .OUT(na1749_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1750_1), .IN8(na1054_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1749_2 ( .OUT(na1749_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1749_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1749_4 ( .OUT(na1749_2_i), .IN1(na1436_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1467_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1749_5 ( .OUT(na1749_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1749_2_i) );
// C_AND////      x98y81     80'h00_0018_00_0000_0888_8811
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1750_1 ( .OUT(na1750_1), .IN1(~na7596_1), .IN2(~na7594_2), .IN3(~na7600_2), .IN4(~na7598_1), .IN5(na7595_1), .IN6(na7597_2),
                      .IN7(na7599_1), .IN8(na7593_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x88y94     80'h00_FE00_80_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1755_4 ( .OUT(na1755_2_i), .IN1(na9954_2), .IN2(~na7601_1), .IN3(na433_2), .IN4(na9228_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1755_5 ( .OUT(na1755_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1755_2_i) );
// C_AND/D///      x89y91     80'h00_FE00_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1758_1 ( .OUT(na1758_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9954_2), .IN6(~na7605_1), .IN7(na9227_2),
                      .IN8(~na452_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1758_2 ( .OUT(na1758_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1758_1_i) );
// C_ORAND/D///      x116y68     80'h00_FE00_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1761_1 ( .OUT(na1761_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7609_1), .IN6(na7610_2), .IN7(1'b0), .IN8(na1762_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1761_2 ( .OUT(na1761_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1761_1_i) );
// C_///AND/      x106y66     80'h00_0060_00_0000_0C08_FF23
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1762_4 ( .OUT(na1762_2), .IN1(1'b1), .IN2(~na435_1), .IN3(na433_2), .IN4(~na452_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x121y72     80'h00_FE00_80_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1764_4 ( .OUT(na1764_2_i), .IN1(na7612_2), .IN2(~na7611_1), .IN3(1'b0), .IN4(na1762_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1764_5 ( .OUT(na1764_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1764_2_i) );
// C_///ORAND/D      x122y74     80'h00_FE00_80_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1766_4 ( .OUT(na1766_2_i), .IN1(na7614_1), .IN2(~na7613_2), .IN3(1'b0), .IN4(na1762_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1766_5 ( .OUT(na1766_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1766_2_i) );
// C_ORAND/D///      x115y69     80'h00_FE00_00_0000_0C88_CBFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1768_1 ( .OUT(na1768_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7616_1), .IN6(~na7615_1), .IN7(1'b0), .IN8(na1762_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1768_2 ( .OUT(na1768_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1768_1_i) );
// C_AND/D//AND/D      x102y72     80'h00_FE00_80_0000_0C88_C38F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1770_1 ( .OUT(na1770_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na7617_1), .IN7(1'b1), .IN8(na1762_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1770_2 ( .OUT(na1770_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1770_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1770_4 ( .OUT(na1770_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na427_2), .IN4(na455_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1770_5 ( .OUT(na1770_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1770_2_i) );
// C_AND/D//AND/D      x103y72     80'h00_FE00_80_0000_0C88_C3AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1774_1 ( .OUT(na1774_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na7623_1), .IN7(1'b1), .IN8(na1762_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1774_2 ( .OUT(na1774_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1774_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1774_4 ( .OUT(na1774_2_i), .IN1(na425_1), .IN2(1'b1), .IN3(na427_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1774_5 ( .OUT(na1774_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1774_2_i) );
// C_AND/D///      x106y76     80'h00_FE00_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1776_1 ( .OUT(na1776_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na7627_1), .IN8(na1762_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1776_2 ( .OUT(na1776_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1776_1_i) );
// C_AND/D///      x88y91     80'h00_FE00_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1780_1 ( .OUT(na1780_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7633_1), .IN6(na435_2), .IN7(na9227_2),
                      .IN8(~na452_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1780_2 ( .OUT(na1780_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1780_1_i) );
// C_AND/D///      x91y91     80'h00_FE00_00_0000_0C88_14FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1783_1 ( .OUT(na1783_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9231_2), .IN6(na435_1), .IN7(~na7637_1),
                      .IN8(~na452_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1783_2 ( .OUT(na1783_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1783_1_i) );
// C_///AND/D      x87y92     80'h00_FE00_80_0000_0C08_FF18
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1786_4 ( .OUT(na1786_2_i), .IN1(na566_1), .IN2(na435_2), .IN3(~na9227_2), .IN4(~na7641_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1786_5 ( .OUT(na1786_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1786_2_i) );
// C_AND/D//AND/D      x86y88     80'h00_FE00_80_0000_0C88_2222
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1792_1 ( .OUT(na1792_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na566_1), .IN6(~na435_1), .IN7(na433_2),
                      .IN8(~na7649_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1792_2 ( .OUT(na1792_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1792_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1792_4 ( .OUT(na1792_2_i), .IN1(na566_1), .IN2(~na435_1), .IN3(na433_1), .IN4(~na7645_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1792_5 ( .OUT(na1792_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1792_2_i) );
// C_///AND/D      x89y92     80'h00_FE00_80_0000_0C08_FF21
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1795_4 ( .OUT(na1795_2_i), .IN1(~na7653_1), .IN2(~na435_1), .IN3(na9265_2), .IN4(~na452_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1795_5 ( .OUT(na1795_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1795_2_i) );
// C_///AND/D      x91y91     80'h00_FE00_80_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1798_4 ( .OUT(na1798_2_i), .IN1(~na7657_1), .IN2(na435_2), .IN3(na9224_2), .IN4(~na9228_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1798_5 ( .OUT(na1798_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1798_2_i) );
// C_///ORAND/D      x98y88     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1801_4 ( .OUT(na1801_2_i), .IN1(~na7661_1), .IN2(na7662_2), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1801_5 ( .OUT(na1801_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1801_2_i) );
// C_MX4b/D///      x93y103     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1803_1 ( .OUT(na1803_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1803_1), .IN6(na1101_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a1803_2 ( .OUT(na1803_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1803_1_i) );
// C_///ORAND/D      x102y90     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1804_4 ( .OUT(na1804_2_i), .IN1(na7664_2), .IN2(~na7663_2), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1804_5 ( .OUT(na1804_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1804_2_i) );
// C_///ORAND/D      x94y97     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1806_4 ( .OUT(na1806_2_i), .IN1(na7666_2), .IN2(~na7665_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1806_5 ( .OUT(na1806_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1806_2_i) );
// C_ORAND/D///      x106y94     80'h00_FE00_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1808_1 ( .OUT(na1808_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7667_1), .IN6(na7668_2), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1808_2 ( .OUT(na1808_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1808_1_i) );
// C_///ORAND/D      x106y95     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1810_4 ( .OUT(na1810_2_i), .IN1(na7670_2), .IN2(~na7669_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1810_5 ( .OUT(na1810_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1810_2_i) );
// C_///ORAND/D      x98y90     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1812_4 ( .OUT(na1812_2_i), .IN1(na7672_1), .IN2(~na7671_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1812_5 ( .OUT(na1812_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1812_2_i) );
// C_ORAND/D///      x94y90     80'h00_FE00_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1814_1 ( .OUT(na1814_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7674_2), .IN6(~na7673_1), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1814_2 ( .OUT(na1814_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1814_1_i) );
// C_///ORAND/D      x100y95     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1816_4 ( .OUT(na1816_2_i), .IN1(~na7675_1), .IN2(na7676_2), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1816_5 ( .OUT(na1816_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1816_2_i) );
// C_ORAND/D///      x96y91     80'h00_FE00_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1818_1 ( .OUT(na1818_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7678_2), .IN6(~na7677_1), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1818_2 ( .OUT(na1818_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1818_1_i) );
// C_ORAND/D///      x104y93     80'h00_FE00_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1820_1 ( .OUT(na1820_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7680_2), .IN6(~na7679_1), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1820_2 ( .OUT(na1820_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1820_1_i) );
// C_///ORAND/D      x106y97     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1822_4 ( .OUT(na1822_2_i), .IN1(na7682_2), .IN2(~na7681_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1822_5 ( .OUT(na1822_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1822_2_i) );
// C_///ORAND/D      x105y94     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1824_4 ( .OUT(na1824_2_i), .IN1(na7684_2), .IN2(~na7683_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1824_5 ( .OUT(na1824_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1824_2_i) );
// C_///ORAND/D      x108y93     80'h00_FE00_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1826_4 ( .OUT(na1826_2_i), .IN1(na7686_2), .IN2(~na7685_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1826_5 ( .OUT(na1826_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1826_2_i) );
// C_MX4b/D///      x123y63     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1828_1 ( .OUT(na1828_1_i), .IN1(na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1828_1), .IN6(na6482_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1828_2 ( .OUT(na1828_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1828_1_i) );
// C_MX4b/D///      x98y99     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1829_1 ( .OUT(na1829_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1829_1),
                      .IN8(na3771_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1829_2 ( .OUT(na1829_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1829_1_i) );
// C_///ORAND/D      x105y93     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1830_4 ( .OUT(na1830_2_i), .IN1(~na7687_1), .IN2(na7688_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1830_5 ( .OUT(na1830_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1830_2_i) );
// C_///ORAND/D      x97y90     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1832_4 ( .OUT(na1832_2_i), .IN1(~na7689_2), .IN2(na7690_2), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1832_5 ( .OUT(na1832_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1832_2_i) );
// C_ORAND/D///      x108y94     80'h00_FE00_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1834_1 ( .OUT(na1834_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7691_2), .IN6(na7692_1), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1834_2 ( .OUT(na1834_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1834_1_i) );
// C_///ORAND/D      x104y93     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1836_4 ( .OUT(na1836_2_i), .IN1(~na7693_2), .IN2(na7694_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1836_5 ( .OUT(na1836_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1836_2_i) );
// C_ORAND/D///      x100y102     80'h00_FE00_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1838_1 ( .OUT(na1838_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7695_2), .IN6(na7696_1), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1838_2 ( .OUT(na1838_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1838_1_i) );
// C_ORAND/D//ORAND/D      x107y76     80'h00_FE00_80_0000_0C88_ADCB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1840_1 ( .OUT(na1840_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7697_2), .IN6(na7698_1), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1840_2 ( .OUT(na1840_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1840_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1840_4 ( .OUT(na1840_2_i), .IN1(na7622_1), .IN2(~na7621_2), .IN3(1'b0), .IN4(na1762_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1840_5 ( .OUT(na1840_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1840_2_i) );
// C_///ORAND/D      x105y95     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1842_4 ( .OUT(na1842_2_i), .IN1(~na7699_1), .IN2(na7700_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1842_5 ( .OUT(na1842_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1842_2_i) );
// C_ORAND/D///      x103y92     80'h00_FE00_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1844_1 ( .OUT(na1844_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7702_1), .IN6(~na7701_2), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1844_2 ( .OUT(na1844_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1844_1_i) );
// C_///ORAND/D      x107y91     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1846_4 ( .OUT(na1846_2_i), .IN1(~na7703_2), .IN2(na7704_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1846_5 ( .OUT(na1846_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1846_2_i) );
// C_///ORAND/D      x101y90     80'h00_FE00_80_0000_0C08_FFAD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1848_4 ( .OUT(na1848_2_i), .IN1(~na7705_2), .IN2(na7706_1), .IN3(na855_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1848_5 ( .OUT(na1848_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1848_2_i) );
// C_ORAND/D///      x101y90     80'h00_FE00_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1850_1 ( .OUT(na1850_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7707_2), .IN6(na7708_2), .IN7(na855_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1850_2 ( .OUT(na1850_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1850_1_i) );
// C_///AND/D      x99y80     80'h00_FE00_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1852_4 ( .OUT(na1852_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na855_1), .IN4(~na7709_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1852_5 ( .OUT(na1852_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1852_2_i) );
// C_MX4b/D///      x95y75     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1854_1 ( .OUT(na1854_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1854_1), .IN6(~na18_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1854_2 ( .OUT(na1854_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1854_1_i) );
// C_MX4b/D///      x95y76     80'h00_FE00_00_0040_0A31_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1855_1 ( .OUT(na1855_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na17_1), .IN6(na1855_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1855_2 ( .OUT(na1855_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1855_1_i) );
// C_AND/D///      x94y97     80'h00_FE00_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1856_1 ( .OUT(na1856_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na7713_1), .IN7(na855_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1856_2 ( .OUT(na1856_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1856_1_i) );
// C_MX4b/D///      x90y63     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1858_1 ( .OUT(na1858_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9534_2), .IN6(na89_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1858_2 ( .OUT(na1858_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1858_1_i) );
// C_AND/D//AND/D      x88y122     80'h00_FE00_80_0000_0C88_F83A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1859_1 ( .OUT(na1859_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na324_1), .IN6(na3892_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1859_2 ( .OUT(na1859_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1859_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1859_4 ( .OUT(na1859_2_i), .IN1(na324_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1859_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1859_5 ( .OUT(na1859_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1859_2_i) );
// C_AND/D///      x97y93     80'h00_FE00_00_0000_0888_1421
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1860_1 ( .OUT(na1860_1_i), .IN1(~na9940_2), .IN2(~na5223_2), .IN3(na3357_1), .IN4(~na3423_1), .IN5(~na3297_2), .IN6(na3600_1),
                      .IN7(~na3292_1), .IN8(~na9812_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1860_2 ( .OUT(na1860_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1860_1_i) );
// C_///AND/D      x104y75     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1861_4 ( .OUT(na1861_2_i), .IN1(na948_1), .IN2(1'b1), .IN3(1'b1), .IN4(na947_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1861_5 ( .OUT(na1861_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1861_2_i) );
// C_MX4b/D///      x105y73     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1863_1 ( .OUT(na1863_1_i), .IN1(1'b1), .IN2(na161_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1863_1), .IN6(na6483_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1863_2 ( .OUT(na1863_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1863_1_i) );
// C_AND/D//AND/D      x80y98     80'h00_F600_80_0000_0C88_F83C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1864_1 ( .OUT(na1864_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3698_2), .IN6(na410_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1864_2 ( .OUT(na1864_1), .CLK(na4116_1), .EN(~na56_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1864_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1864_4 ( .OUT(na1864_2_i), .IN1(1'b1), .IN2(na410_1), .IN3(1'b1), .IN4(~na1864_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1864_5 ( .OUT(na1864_2), .CLK(na4116_1), .EN(~na56_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1864_2_i) );
// C_AND////      x98y72     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1865_1 ( .OUT(na1865_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9947_2), .IN6(1'b1), .IN7(1'b1), .IN8(na73_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x101y69     80'h00_0018_00_0000_0C88_63FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1866_1 ( .OUT(na1866_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na36_2), .IN7(na6684_2), .IN8(~na6673_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x101y101     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1867_1 ( .OUT(na1867_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1867_1), .IN6(na1091_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1867_2 ( .OUT(na1867_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1867_1_i) );
// C_MX4b/D///      x115y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1868_1 ( .OUT(na1868_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1868_1), .IN6(na1103_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1868_2 ( .OUT(na1868_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1868_1_i) );
// C_MX4b/D///      x117y89     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1869_1 ( .OUT(na1869_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1869_1), .IN6(na1101_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1869_2 ( .OUT(na1869_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1869_1_i) );
// C_MX4b/D///      x95y93     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1870_1 ( .OUT(na1870_1_i), .IN1(na954_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1870_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1870_2 ( .OUT(na1870_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1870_1_i) );
// C_MX2a////      x84y79     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1872_1 ( .OUT(na1872_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1065_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1067_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x92y89     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1875_1 ( .OUT(na1875_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na913_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na915_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y87     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1877_1 ( .OUT(na1877_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1337_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1339_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y91     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1879_1 ( .OUT(na1879_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1061_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1063_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x93y62     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1880_4 ( .OUT(na1880_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1881_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1880_5 ( .OUT(na1880_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1880_2_i) );
// C_MX2a////      x92y77     80'h00_0018_00_0040_0CAA_8F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1881_1 ( .OUT(na1881_1), .IN1(1'b0), .IN2(~na1880_2), .IN3(1'b0), .IN4(~na159_1), .IN5(1'b1), .IN6(1'b1), .IN7(na436_1),
                      .IN8(na1882_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y76     80'h00_0018_00_0000_0C88_82FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1882_1 ( .OUT(na1882_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(~na435_1), .IN7(na433_1), .IN8(na9223_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x119y93     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1883_1 ( .OUT(na1883_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1883_1), .IN6(na1105_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1883_2 ( .OUT(na1883_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1883_1_i) );
// C_MX4b/D///      x101y72     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1885_1 ( .OUT(na1885_1_i), .IN1(1'b1), .IN2(na161_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9536_2),
                      .IN8(na6478_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1885_2 ( .OUT(na1885_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1885_1_i) );
// C_AND/D///      x84y83     80'h00_FE00_00_0000_0888_38F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1886_1 ( .OUT(na1886_1_i), .IN1(na428_1), .IN2(na435_1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(na942_1), .IN7(1'b1),
                      .IN8(~na452_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1886_2 ( .OUT(na1886_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1886_1_i) );
// C_AND/D//AND/D      x49y120     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1888_1 ( .OUT(na1888_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3826_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1888_2 ( .OUT(na1888_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1888_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1888_4 ( .OUT(na1888_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(na3826_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1888_5 ( .OUT(na1888_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1888_2_i) );
// C_MX4b/D///      x119y79     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1889_1 ( .OUT(na1889_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na9537_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1889_2 ( .OUT(na1889_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1889_1_i) );
// C_MX4b/D///      x110y81     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1891_1 ( .OUT(na1891_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1891_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1891_2 ( .OUT(na1891_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1891_1_i) );
// C_MX4b/D///      x112y79     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1892_1 ( .OUT(na1892_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1892_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1892_2 ( .OUT(na1892_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1892_1_i) );
// C_MX4b/D///      x116y64     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1893_1 ( .OUT(na1893_1_i), .IN1(~na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na1893_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1893_2 ( .OUT(na1893_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1893_1_i) );
// C_MX4b/D///      x120y66     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1894_1 ( .OUT(na1894_1_i), .IN1(~na876_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na1894_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1894_2 ( .OUT(na1894_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1894_1_i) );
// C_///AND/D      x110y71     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1895_4 ( .OUT(na1895_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1896_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1895_5 ( .OUT(na1895_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1895_2_i) );
// C_MX2a////      x106y79     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1896_1 ( .OUT(na1896_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1895_2), .IN4(~na159_1), .IN5(na853_2), .IN6(na873_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x95y105     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1897_1 ( .OUT(na1897_1_i), .IN1(na569_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1897_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1897_2 ( .OUT(na1897_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1897_1_i) );
// C_MX4b/D///      x95y112     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1898_1 ( .OUT(na1898_1_i), .IN1(~na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na5185_1), .IN6(na1898_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1898_2 ( .OUT(na1898_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1898_1_i) );
// C_MX4b/D///      x95y111     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1899_1 ( .OUT(na1899_1_i), .IN1(na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1899_1), .IN6(na5181_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1899_2 ( .OUT(na1899_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1899_1_i) );
// C_AND/D///      x103y95     80'h00_FE00_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1900_1 ( .OUT(na1900_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1275_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1900_2 ( .OUT(na1900_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1900_1_i) );
// C_MX4b/D///      x111y103     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1901_1 ( .OUT(na1901_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2667_1), .IN6(~na1902_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1901_2 ( .OUT(na1901_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1901_1_i) );
// C_MX2b////      x105y106     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1902_1 ( .OUT(na1902_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1275_1), .IN4(1'b1), .IN5(~na4012_1), .IN6(1'b0), .IN7(~na9461_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x97y101     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1903_1 ( .OUT(na1903_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3750_2),
                      .IN8(na9540_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1903_2 ( .OUT(na1903_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1903_1_i) );
// C_ORAND*////D      x88y71     80'h00_FE18_00_0000_0788_37BC
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1904_1 ( .OUT(na1904_1), .IN1(1'b0), .IN2(na1917_1), .IN3(na1905_1), .IN4(~na1921_1), .IN5(~na2947_1), .IN6(~na9542_2), .IN7(1'b0),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1904_5 ( .OUT(na1904_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1904_1) );
// C_AND////      x94y83     80'h00_0018_00_0000_0888_2128
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1905_1 ( .OUT(na1905_1), .IN1(na1915_1), .IN2(na1907_1), .IN3(na1914_1), .IN4(~na3143_1), .IN5(~na1915_2), .IN6(~na1479_1),
                      .IN7(na1914_2), .IN8(~na3198_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y88     80'h00_0018_00_0000_0888_3128
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1907_1 ( .OUT(na1907_1), .IN1(na1911_2), .IN2(na1909_1), .IN3(na1910_2), .IN4(~na1792_1), .IN5(~na1783_1), .IN6(~na1786_2),
                      .IN7(1'b1), .IN8(~na1792_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y86     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1909_1 ( .OUT(na1909_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1798_2), .IN6(~na1795_2), .IN7(~na3554_1),
                      .IN8(~na1590_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y91     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1910_4 ( .OUT(na1910_2), .IN1(~na1758_1), .IN2(~na1545_2), .IN3(~na1780_1), .IN4(~na1755_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y87     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1911_4 ( .OUT(na1911_2), .IN1(~na1040_1), .IN2(~na1542_1), .IN3(~na1538_2), .IN4(~na1475_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y85     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1914_1 ( .OUT(na1914_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1749_2), .IN6(~na1683_2), .IN7(~na1886_1),
                      .IN8(~na3145_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1914_4 ( .OUT(na1914_2), .IN1(~na1749_1), .IN2(~na1683_1), .IN3(~na3149_1), .IN4(~na3559_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y71     80'h00_0078_00_0000_0C88_11AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1915_1 ( .OUT(na1915_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2835_2), .IN6(~na1568_2), .IN7(~na1856_1),
                      .IN8(~na1776_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1915_4 ( .OUT(na1915_2), .IN1(na2835_1), .IN2(1'b1), .IN3(na6455_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y60     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1917_1 ( .OUT(na1917_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1918_1), .IN8(na1920_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y49     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1918_1 ( .OUT(na1918_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9366_2), .IN6(~na7723_1), .IN7(~na977_2),
                      .IN8(~na9950_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x82y58     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1920_4 ( .OUT(na1920_2), .IN1(~na9368_2), .IN2(~na9956_2), .IN3(~na977_1), .IN4(~na10040_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x88y70     80'h00_0078_00_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1921_1 ( .OUT(na1921_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na979_1), .IN7(na1113_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1921_4 ( .OUT(na1921_2), .IN1(na214_2), .IN2(1'b1), .IN3(na978_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x82y65     80'h00_FE18_00_0000_0EEE_E3E0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1922_1 ( .OUT(na1922_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1930_2), .IN4(na1929_1), .IN5(1'b0), .IN6(~na7730_1), .IN7(na1930_1),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1922_5 ( .OUT(na1922_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1922_1) );
// C_///AND/      x106y68     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1927_4 ( .OUT(na1927_2), .IN1(~na1473_2), .IN2(~na1852_2), .IN3(~na1564_2), .IN4(~na1535_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y56     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1929_1 ( .OUT(na1929_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7732_1), .IN7(na977_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x86y71     80'h00_0078_00_0000_0C88_AACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1930_1 ( .OUT(na1930_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7733_1), .IN6(1'b1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1930_4 ( .OUT(na1930_2), .IN1(1'b1), .IN2(na7727_1), .IN3(1'b1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y66     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1931_1 ( .OUT(na1931_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6386_1), .IN6(~na6385_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x84y69     80'h00_FE18_00_0000_0EEE_EAA3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1932_1 ( .OUT(na1932_1), .IN1(1'b0), .IN2(~na7738_1), .IN3(na1940_1), .IN4(1'b0), .IN5(na1939_1), .IN6(1'b0), .IN7(na1940_2),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1932_5 ( .OUT(na1932_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1932_1) );
// C_AND////      x108y70     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1937_1 ( .OUT(na1937_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1562_2), .IN6(~na1850_1), .IN7(~na1470_2),
                      .IN8(~na1532_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y53     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1939_1 ( .OUT(na1939_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na977_2), .IN8(na7740_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x86y69     80'h00_0078_00_0000_0C88_8FCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1940_1 ( .OUT(na1940_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na977_1), .IN8(na7741_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1940_4 ( .OUT(na1940_2), .IN1(1'b1), .IN2(na7735_1), .IN3(1'b1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y61     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1941_1 ( .OUT(na1941_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6388_1), .IN6(~na6387_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x84y68     80'h00_FE18_00_0000_0EEE_CA3E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1942_1 ( .OUT(na1942_1), .IN1(na1949_2), .IN2(na1944_2), .IN3(1'b0), .IN4(~na7743_2), .IN5(na1949_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1942_5 ( .OUT(na1942_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1942_1) );
// C_///AND/      x93y66     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1944_4 ( .OUT(na1944_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_2), .IN4(na7745_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x85y69     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1949_1 ( .OUT(na1949_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7749_1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1949_4 ( .OUT(na1949_2), .IN1(na9541_2), .IN2(1'b1), .IN3(1'b1), .IN4(na7746_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y61     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1950_1 ( .OUT(na1950_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6390_1), .IN6(~na6389_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x83y68     80'h00_FE18_00_0000_0EEE_CAAB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1951_1 ( .OUT(na1951_1), .IN1(na1958_2), .IN2(~na7751_2), .IN3(na1953_2), .IN4(1'b0), .IN5(na1958_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1951_5 ( .OUT(na1951_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1951_1) );
// C_///AND/      x80y61     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1953_4 ( .OUT(na1953_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_2), .IN4(na7753_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x85y67     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1958_1 ( .OUT(na1958_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7757_1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1958_4 ( .OUT(na1958_2), .IN1(na9541_2), .IN2(1'b1), .IN3(1'b1), .IN4(na7754_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y58     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1959_1 ( .OUT(na1959_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6392_1), .IN6(~na6391_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x81y69     80'h00_FE18_00_0000_0EEE_CBAA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1960_1 ( .OUT(na1960_1), .IN1(na1967_2), .IN2(1'b0), .IN3(na1962_2), .IN4(1'b0), .IN5(na1967_1), .IN6(~na7759_2), .IN7(1'b0),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1960_5 ( .OUT(na1960_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1960_1) );
// C_///AND/      x84y73     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1962_4 ( .OUT(na1962_2), .IN1(1'b1), .IN2(na7761_1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x83y67     80'h00_0078_00_0000_0C88_8FCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1967_1 ( .OUT(na1967_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na977_1), .IN8(na7765_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1967_4 ( .OUT(na1967_2), .IN1(na7762_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y62     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1968_1 ( .OUT(na1968_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6394_1), .IN6(~na6393_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x83y72     80'h00_FE18_00_0000_0EEE_E0BA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1969_1 ( .OUT(na1969_1), .IN1(na1971_2), .IN2(1'b0), .IN3(na1976_2), .IN4(~na7767_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1976_1),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1969_5 ( .OUT(na1969_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1969_1) );
// C_///AND/      x83y75     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1971_4 ( .OUT(na1971_2), .IN1(na7769_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x86y67     80'h00_0078_00_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1976_1 ( .OUT(na1976_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9366_2), .IN6(1'b1), .IN7(na7773_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1976_4 ( .OUT(na1976_2), .IN1(1'b1), .IN2(1'b1), .IN3(na7770_1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x62y49     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1977_1 ( .OUT(na1977_1), .IN1(1'b1), .IN2(1'b1), .IN3(na90_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na6395_1), .IN7(1'b0), .IN8(~na6396_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x83y65     80'h00_FE18_00_0000_0EEE_E0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1978_1 ( .OUT(na1978_1), .IN1(1'b0), .IN2(na1980_1), .IN3(na1981_1), .IN4(na7774_2), .IN5(1'b0), .IN6(1'b0), .IN7(na9188_2),
                      .IN8(na7774_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1978_5 ( .OUT(na1978_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1978_1) );
// C_AND////      x93y74     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1980_1 ( .OUT(na1980_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na2938_1), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y59     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1981_1 ( .OUT(na1981_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9367_2), .IN6(1'b1), .IN7(na7775_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x78y57     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1982_1 ( .OUT(na1982_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6398_1), .IN6(~na6397_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y64     80'h00_0018_00_0000_0888_5123
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1984_1 ( .OUT(na1984_1), .IN1(1'b1), .IN2(~na1840_1), .IN3(na1986_2), .IN4(~na1435_1), .IN5(~na1741_1), .IN6(~na1840_2),
                      .IN7(~na1669_2), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y83     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1986_4 ( .OUT(na1986_2), .IN1(~na1597_1), .IN2(~na1509_1), .IN3(~na1548_2), .IN4(~na1571_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x84y66     80'h00_FE18_00_0000_0EEE_E3AA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1987_1 ( .OUT(na1987_1), .IN1(na7780_1), .IN2(1'b0), .IN3(na1990_2), .IN4(1'b0), .IN5(1'b0), .IN6(~na7778_2), .IN7(na1990_1),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1987_5 ( .OUT(na1987_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1987_1) );
// C_AND///AND/      x82y61     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1990_1 ( .OUT(na1990_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7781_1), .IN7(na977_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1990_4 ( .OUT(na1990_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_1), .IN4(na7782_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y74     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1991_4 ( .OUT(na1991_2), .IN1(~na1667_1), .IN2(~na1739_2), .IN3(~na1506_2), .IN4(~na1838_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y66     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1993_1 ( .OUT(na1993_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6399_1), .IN8(na6400_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x82y66     80'h00_FE18_00_0000_0EEE_BACA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1994_1 ( .OUT(na1994_1), .IN1(na1997_2), .IN2(1'b0), .IN3(1'b0), .IN4(na7786_1), .IN5(na1997_1), .IN6(1'b0), .IN7(na9188_2),
                      .IN8(~na7784_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1994_5 ( .OUT(na1994_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1994_1) );
// C_AND///AND/      x83y61     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1997_1 ( .OUT(na1997_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7787_1), .IN7(na977_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1997_4 ( .OUT(na1997_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_1), .IN4(na7788_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y89     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1998_1 ( .OUT(na1998_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1420_2), .IN6(~na1737_1), .IN7(~na1836_2),
                      .IN8(~na1665_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y64     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2000_1 ( .OUT(na2000_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6401_1), .IN6(na6402_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x82y70     80'h00_FE18_00_0000_0EEE_D0EC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2001_1 ( .OUT(na2001_1), .IN1(1'b0), .IN2(na7792_1), .IN3(na9548_2), .IN4(na2004_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na7790_1),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2001_5 ( .OUT(na2001_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2001_1) );
// C_AND///AND/      x80y60     80'h00_0078_00_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2004_1 ( .OUT(na2004_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7793_1), .IN7(na977_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2004_4 ( .OUT(na2004_2), .IN1(na7794_1), .IN2(1'b1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x110y68     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2005_4 ( .OUT(na2005_2), .IN1(~na1431_2), .IN2(~na1735_1), .IN3(~na1663_1), .IN4(~na1834_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y63     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2007_1 ( .OUT(na2007_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6404_1), .IN8(na6403_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x77y68     80'h00_FE18_00_0000_0EEE_DACA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2008_1 ( .OUT(na2008_1), .IN1(na2011_2), .IN2(1'b0), .IN3(1'b0), .IN4(na7798_1), .IN5(na2011_1), .IN6(1'b0), .IN7(~na7796_2),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2008_5 ( .OUT(na2008_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2008_1) );
// C_AND///AND/      x77y63     80'h00_0078_00_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2011_1 ( .OUT(na2011_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na977_2), .IN8(na7799_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2011_4 ( .OUT(na2011_2), .IN1(na7800_1), .IN2(1'b1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y70     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2012_4 ( .OUT(na2012_2), .IN1(~na1733_2), .IN2(~na1832_2), .IN3(~na1490_1), .IN4(~na1659_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y65     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2014_1 ( .OUT(na2014_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6406_1), .IN6(na6405_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x80y64     80'h00_FE18_00_0000_0EEE_CC3E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2015_1 ( .OUT(na2015_1), .IN1(na7804_1), .IN2(na2018_2), .IN3(1'b0), .IN4(~na7802_2), .IN5(1'b0), .IN6(na2018_1), .IN7(1'b0),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2015_5 ( .OUT(na2015_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2015_1) );
// C_AND///AND/      x81y64     80'h00_0078_00_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2018_1 ( .OUT(na2018_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na977_2), .IN8(na7805_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2018_4 ( .OUT(na2018_2), .IN1(1'b1), .IN2(na7806_1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y69     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2019_4 ( .OUT(na2019_2), .IN1(~na1830_2), .IN2(~na1731_2), .IN3(~na1661_2), .IN4(~na1488_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y64     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2021_1 ( .OUT(na2021_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6407_1), .IN6(na6408_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x86y68     80'h00_FE18_00_0000_0EEE_E5E0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2022_1 ( .OUT(na2022_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2025_2), .IN4(na7810_1), .IN5(~na7808_2), .IN6(1'b0), .IN7(na2025_1),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2022_5 ( .OUT(na2022_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2022_1) );
// C_AND///AND/      x84y63     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2025_1 ( .OUT(na2025_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7811_1), .IN6(1'b1), .IN7(na977_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2025_4 ( .OUT(na2025_2), .IN1(na7812_1), .IN2(1'b1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y74     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2026_1 ( .OUT(na2026_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1486_1), .IN6(~na1390_2), .IN7(~na851_2),
                      .IN8(~na1654_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y62     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2028_1 ( .OUT(na2028_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6410_1), .IN8(na6409_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x86y72     80'h00_FE18_00_0000_0EEE_CBCA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2029_1 ( .OUT(na2029_1), .IN1(na2032_2), .IN2(1'b0), .IN3(1'b0), .IN4(na7816_2), .IN5(na2032_1), .IN6(~na7814_2), .IN7(1'b0),
                      .IN8(na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2029_5 ( .OUT(na2029_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2029_1) );
// C_AND///AND/      x81y61     80'h00_0078_00_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2032_1 ( .OUT(na2032_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7817_1), .IN6(1'b1), .IN7(na977_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2032_4 ( .OUT(na2032_2), .IN1(1'b1), .IN2(na7818_1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y72     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2033_1 ( .OUT(na2033_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1484_2), .IN6(~na1651_1), .IN7(~na1401_2),
                      .IN8(~na861_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y65     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2035_1 ( .OUT(na2035_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6412_1), .IN6(na6411_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////D      x83y64     80'h00_FE18_00_0000_0EEE_BCCC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2036_1 ( .OUT(na2036_1), .IN1(1'b0), .IN2(na2039_2), .IN3(1'b0), .IN4(na7822_1), .IN5(1'b0), .IN6(na2039_1), .IN7(na9188_2),
                      .IN8(~na7820_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2036_5 ( .OUT(na2036_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2036_1) );
// C_AND///AND/      x87y60     80'h00_0078_00_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2039_1 ( .OUT(na2039_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7823_1), .IN6(1'b1), .IN7(na977_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2039_4 ( .OUT(na2039_2), .IN1(na7824_1), .IN2(1'b1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y73     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2040_1 ( .OUT(na2040_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1724_1), .IN6(~na1649_2), .IN7(~na1482_1),
                      .IN8(~na884_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y63     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2042_1 ( .OUT(na2042_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6413_1), .IN8(na6414_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x85y66     80'h00_FE18_00_0000_0788_3551
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2043_1 ( .OUT(na2043_1), .IN1(~na2045_2), .IN2(~na2048_1), .IN3(~na2046_1), .IN4(1'b1), .IN5(~na2045_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2043_5 ( .OUT(na2043_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2043_1) );
// C_AND///AND/      x93y67     80'h00_0078_00_0000_0C88_A88F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2045_1 ( .OUT(na2045_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na891_1), .IN6(na9185_2), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2045_4 ( .OUT(na2045_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_2), .IN4(na7828_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y61     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2046_1 ( .OUT(na2046_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7825_1), .IN6(1'b1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y62     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2047_1 ( .OUT(na2047_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6415_1), .IN6(~na6416_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y66     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2048_1 ( .OUT(na2048_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9541_2), .IN6(1'b1), .IN7(1'b1), .IN8(na7826_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x85y72     80'h00_FE18_00_0000_0788_3153
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2050_1 ( .OUT(na2050_1), .IN1(1'b1), .IN2(~na2052_2), .IN3(~na2055_1), .IN4(1'b1), .IN5(~na2053_2), .IN6(~na2052_1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2050_5 ( .OUT(na2050_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2050_1) );
// C_AND///AND/      x93y68     80'h00_0078_00_0000_0C88_A8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2052_1 ( .OUT(na2052_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na1885_1), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2052_4 ( .OUT(na2052_2), .IN1(na7832_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y59     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2053_4 ( .OUT(na2053_2), .IN1(na9367_2), .IN2(1'b1), .IN3(na7829_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y60     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2054_1 ( .OUT(na2054_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6418_1), .IN6(~na6417_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y73     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2055_1 ( .OUT(na2055_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9541_2), .IN6(1'b1), .IN7(1'b1), .IN8(na7830_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x81y68     80'h00_FE18_00_0000_0788_3551
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2057_1 ( .OUT(na2057_1), .IN1(~na2059_2), .IN2(~na2060_2), .IN3(~na2062_1), .IN4(1'b1), .IN5(~na2059_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2057_5 ( .OUT(na2057_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2057_1) );
// C_AND///AND/      x91y67     80'h00_0078_00_0000_0C88_8AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2059_1 ( .OUT(na2059_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na160_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2059_4 ( .OUT(na2059_2), .IN1(na7836_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y60     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2060_4 ( .OUT(na2060_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_1), .IN4(na7833_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y55     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2061_1 ( .OUT(na2061_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6419_1), .IN6(~na6420_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y73     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2062_1 ( .OUT(na2062_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7834_1), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x84y70     80'h00_FE18_00_0000_0788_3551
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2064_1 ( .OUT(na2064_1), .IN1(~na2066_2), .IN2(~na2067_2), .IN3(~na2069_2), .IN4(1'b1), .IN5(~na2066_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2064_5 ( .OUT(na2064_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2064_1) );
// C_AND///AND/      x85y65     80'h00_0078_00_0000_0C88_A8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2066_1 ( .OUT(na2066_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na164_1), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2066_4 ( .OUT(na2066_2), .IN1(na9368_2), .IN2(1'b1), .IN3(na7840_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y58     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2067_4 ( .OUT(na2067_2), .IN1(1'b1), .IN2(na7837_1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y59     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2068_1 ( .OUT(na2068_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6421_1), .IN6(~na6422_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y73     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2069_4 ( .OUT(na2069_2), .IN1(1'b1), .IN2(na7838_2), .IN3(1'b1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x79y68     80'h00_FE18_00_0000_0788_3153
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2071_1 ( .OUT(na2071_1), .IN1(1'b1), .IN2(~na2073_2), .IN3(~na2074_1), .IN4(1'b1), .IN5(~na2076_2), .IN6(~na2073_1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2071_5 ( .OUT(na2071_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2071_1) );
// C_AND///AND/      x87y68     80'h00_0078_00_0000_0C88_8AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2073_1 ( .OUT(na2073_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2073_4 ( .OUT(na2073_2), .IN1(na7844_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y63     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2074_1 ( .OUT(na2074_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na977_1), .IN8(na7841_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y60     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2075_1 ( .OUT(na2075_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na6424_1), .IN8(~na6423_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y71     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2076_4 ( .OUT(na2076_2), .IN1(1'b1), .IN2(1'b1), .IN3(na7842_1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x80y74     80'h00_FE18_00_0000_0788_1F15
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2078_1 ( .OUT(na2078_1), .IN1(~na2081_1), .IN2(1'b1), .IN3(~na2083_1), .IN4(~na2080_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na9188_2),
                      .IN8(~na2080_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2078_5 ( .OUT(na2078_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2078_1) );
// C_AND///AND/      x94y66     80'h00_0078_00_0000_0C88_8AAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2080_1 ( .OUT(na2080_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na166_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2080_4 ( .OUT(na2080_2), .IN1(1'b1), .IN2(na7848_1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y59     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2081_1 ( .OUT(na2081_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7845_1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y60     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2082_1 ( .OUT(na2082_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6426_1), .IN6(~na6425_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y79     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2083_1 ( .OUT(na2083_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7846_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x89y68     80'h00_FE18_00_0000_0788_131F
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2085_1 ( .OUT(na2085_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na2087_2), .IN4(~na2090_2), .IN5(1'b1), .IN6(~na2088_2), .IN7(~na2087_1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2085_5 ( .OUT(na2085_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2085_1) );
// C_AND///AND/      x98y67     80'h00_0078_00_0000_0C88_A88F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2087_1 ( .OUT(na2087_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1863_1), .IN6(na9185_2), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2087_4 ( .OUT(na2087_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_2), .IN4(na7852_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y58     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2088_4 ( .OUT(na2088_2), .IN1(na7849_1), .IN2(1'b1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y55     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2089_1 ( .OUT(na2089_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6427_1), .IN6(~na6428_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y56     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2090_4 ( .OUT(na2090_2), .IN1(na7850_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x85y68     80'h00_FE18_00_0000_0788_3351
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2092_1 ( .OUT(na2092_1), .IN1(~na2097_1), .IN2(~na2094_2), .IN3(~na2095_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2094_1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2092_5 ( .OUT(na2092_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2092_1) );
// C_AND///AND/      x81y60     80'h00_0078_00_0000_0C88_A8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2094_1 ( .OUT(na2094_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na167_1), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2094_4 ( .OUT(na2094_2), .IN1(na9368_2), .IN2(1'b1), .IN3(na7856_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y59     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2095_1 ( .OUT(na2095_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7853_1), .IN6(1'b1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y59     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2096_1 ( .OUT(na2096_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6429_1), .IN6(~na6430_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x103y55     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2097_1 ( .OUT(na2097_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7854_1), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x80y62     80'h00_FE18_00_0000_0788_3351
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2099_1 ( .OUT(na2099_1), .IN1(~na2102_1), .IN2(~na2101_2), .IN3(~na2104_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na2101_1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2099_5 ( .OUT(na2099_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2099_1) );
// C_AND///AND/      x85y64     80'h00_0078_00_0000_0C88_8AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2101_1 ( .OUT(na2101_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na1623_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2101_4 ( .OUT(na2101_2), .IN1(na7860_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y63     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2102_1 ( .OUT(na2102_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7857_1), .IN6(1'b1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y58     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2103_1 ( .OUT(na2103_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6432_1), .IN6(~na6431_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x86y73     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2104_4 ( .OUT(na2104_2), .IN1(na7858_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1921_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x88y62     80'h00_FE18_00_0000_0788_1F51
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2106_1 ( .OUT(na2106_1), .IN1(~na2109_1), .IN2(~na2111_1), .IN3(~na2108_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2108_1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2106_5 ( .OUT(na2106_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2106_1) );
// C_AND///AND/      x94y65     80'h00_0078_00_0000_0C88_A8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2108_1 ( .OUT(na2108_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na267_1), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2108_4 ( .OUT(na2108_2), .IN1(na7864_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y65     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2109_1 ( .OUT(na2109_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na977_1), .IN8(na7861_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y60     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2110_1 ( .OUT(na2110_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6433_1), .IN6(~na6434_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y58     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2111_1 ( .OUT(na2111_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7862_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x84y72     80'h00_FE18_00_0000_0788_151F
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2113_1 ( .OUT(na2113_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na2115_2), .IN4(~na2118_1), .IN5(~na2116_1), .IN6(1'b1), .IN7(~na2115_1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2113_5 ( .OUT(na2113_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2113_1) );
// C_AND///AND/      x88y67     80'h00_0078_00_0000_0C88_8AAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2115_1 ( .OUT(na2115_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na3185_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2115_4 ( .OUT(na2115_2), .IN1(1'b1), .IN2(na7868_1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y63     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2116_1 ( .OUT(na2116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7865_1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y59     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2117_1 ( .OUT(na2117_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6436_1), .IN6(~na6435_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y60     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2118_1 ( .OUT(na2118_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na7866_1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x82y68     80'h00_FE18_00_0000_0788_3313
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2120_1 ( .OUT(na2120_1), .IN1(1'b1), .IN2(~na2122_2), .IN3(~na2123_2), .IN4(~na2125_1), .IN5(1'b1), .IN6(~na2122_1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2120_5 ( .OUT(na2120_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2120_1) );
// C_AND///AND/      x91y66     80'h00_0078_00_0000_0C88_A88F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2122_1 ( .OUT(na2122_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na3177_1), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2122_4 ( .OUT(na2122_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_2), .IN4(na7872_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y61     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2123_4 ( .OUT(na2123_2), .IN1(1'b1), .IN2(na7869_1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y55     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2124_1 ( .OUT(na2124_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na6437_1), .IN8(~na6438_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y58     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2125_1 ( .OUT(na2125_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7870_2), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x82y60     80'h00_FE18_00_0000_0788_3351
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2127_1 ( .OUT(na2127_1), .IN1(~na2132_1), .IN2(~na2129_2), .IN3(~na2130_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na2129_1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2127_5 ( .OUT(na2127_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2127_1) );
// C_AND///AND/      x89y64     80'h00_0078_00_0000_0C88_8AAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2129_1 ( .OUT(na2129_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na3164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2129_4 ( .OUT(na2129_2), .IN1(1'b1), .IN2(na7876_1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y67     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2130_4 ( .OUT(na2130_2), .IN1(1'b1), .IN2(na7873_1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y56     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2131_1 ( .OUT(na2131_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6440_1), .IN6(~na6439_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y55     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2132_1 ( .OUT(na2132_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7874_2), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x80y72     80'h00_FE18_00_0000_0788_1553
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2134_1 ( .OUT(na2134_1), .IN1(1'b1), .IN2(~na9561_2), .IN3(~na2139_1), .IN4(1'b1), .IN5(~na2137_2), .IN6(1'b1), .IN7(~na2136_1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2134_5 ( .OUT(na2134_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2134_1) );
// C_AND///AND/      x90y61     80'h00_0078_00_0000_0C88_8AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2136_1 ( .OUT(na2136_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na3163_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2136_4 ( .OUT(na2136_2), .IN1(na7880_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y65     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2137_4 ( .OUT(na2137_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_1), .IN4(na7877_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y54     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2138_1 ( .OUT(na2138_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na6441_1), .IN8(~na6442_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y59     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2139_1 ( .OUT(na2139_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7878_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x84y60     80'h00_FE18_00_0000_0788_1555
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2141_1 ( .OUT(na2141_1), .IN1(~na9563_2), .IN2(1'b1), .IN3(~na2144_1), .IN4(1'b1), .IN5(~na2146_1), .IN6(1'b1), .IN7(~na2143_1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2141_5 ( .OUT(na2141_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2141_1) );
// C_AND///AND/      x90y65     80'h00_0078_00_0000_0C88_8AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2143_1 ( .OUT(na2143_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(1'b1), .IN7(na978_1), .IN8(na3154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2143_4 ( .OUT(na2143_2), .IN1(na7884_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y57     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2144_1 ( .OUT(na2144_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7881_1), .IN7(na977_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y53     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2145_1 ( .OUT(na2145_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6444_1), .IN6(~na6443_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y57     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2146_1 ( .OUT(na2146_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na7882_2), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x80y68     80'h00_FE18_00_0000_0788_3331
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2148_1 ( .OUT(na2148_1), .IN1(~na2153_1), .IN2(~na2150_2), .IN3(1'b1), .IN4(~na2151_2), .IN5(1'b1), .IN6(~na2150_1), .IN7(1'b1),
                      .IN8(~na228_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2148_5 ( .OUT(na2148_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2148_1) );
// C_AND///AND/      x91y64     80'h00_0078_00_0000_0C88_A88F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2150_1 ( .OUT(na2150_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na3065_1), .IN7(na978_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2150_4 ( .OUT(na2150_2), .IN1(1'b1), .IN2(1'b1), .IN3(na977_2), .IN4(na7888_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x74y68     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2151_4 ( .OUT(na2151_2), .IN1(na7885_1), .IN2(1'b1), .IN3(na977_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y57     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2152_1 ( .OUT(na2152_1), .IN1(1'b1), .IN2(~na9167_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6446_1), .IN6(~na6445_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x109y57     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2153_1 ( .OUT(na2153_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7886_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x84y92     80'h00_FE00_80_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2155_4 ( .OUT(na2155_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4853_2), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2155_5 ( .OUT(na2155_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2155_2_i) );
// C_MX4b/D///      x121y79     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2156_1 ( .OUT(na2156_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2156_1), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2156_2 ( .OUT(na2156_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2156_1_i) );
// C_MX4b/D///      x100y101     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2157_1 ( .OUT(na2157_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2157_1),
                      .IN8(na3767_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2157_2 ( .OUT(na2157_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2157_1_i) );
// C_AND/D//AND/D      x52y110     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2158_1 ( .OUT(na2158_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3831_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2158_2 ( .OUT(na2158_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2158_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2158_4 ( .OUT(na2158_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3831_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2158_5 ( .OUT(na2158_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2158_2_i) );
// C_MX4b/D///      x105y119     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2159_1 ( .OUT(na2159_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1104_1), .IN6(~na2160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2159_2 ( .OUT(na2159_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2159_1_i) );
// C_MX2b////      x107y108     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2160_1 ( .OUT(na2160_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1275_1), .IN4(1'b1), .IN5(~na4007_2), .IN6(1'b0), .IN7(~na9457_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x105y120     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2161_1 ( .OUT(na2161_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1102_1), .IN6(~na2162_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2161_2 ( .OUT(na2161_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2161_1_i) );
// C_MX2b////      x109y106     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2162_1 ( .OUT(na2162_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1275_1), .IN4(1'b1), .IN5(~na4007_1), .IN6(1'b0), .IN7(~na9455_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x116y65     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2163_1 ( .OUT(na2163_1_i), .IN1(na1728_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2163_1),
                      .IN8(na2164_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2163_2 ( .OUT(na2163_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2163_1_i) );
// C_///AND/      x118y58     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2164_4 ( .OUT(na2164_2), .IN1(~na1730_1), .IN2(1'b1), .IN3(na3885_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x99y104     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2165_1 ( .OUT(na2165_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1139_1), .IN6(na2165_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2165_2 ( .OUT(na2165_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2165_1_i) );
// C_MX4b/D///      x102y122     80'h00_FE00_00_0040_0A31_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2166_1 ( .OUT(na2166_1_i), .IN1(~na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na2167_1), .IN6(na2668_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2166_2 ( .OUT(na2166_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2166_1_i) );
// C_MX2b////      x105y103     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2167_1 ( .OUT(na2167_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1275_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na4005_2), .IN7(1'b0), .IN8(~na1205_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x120y80     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2168_1 ( .OUT(na2168_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9564_2), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2168_2 ( .OUT(na2168_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2168_1_i) );
// C_MX4b/D///      x107y101     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2170_1 ( .OUT(na2170_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2170_1), .IN6(na1073_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2170_2 ( .OUT(na2170_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2170_1_i) );
// C_MX2a/D///      x50y120     80'h00_FE00_00_0040_0C8C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2171_1 ( .OUT(na2171_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na9566_2), .IN4(~na527_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2171_2 ( .OUT(na2171_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2171_1_i) );
// C_AND///AND/      x45y118     80'h00_0078_00_0000_0C88_8F8C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2172_1 ( .OUT(na2172_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na359_2), .IN8(na2171_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2172_4 ( .OUT(na2172_2), .IN1(1'b1), .IN2(na504_1), .IN3(na359_1), .IN4(na3324_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x57y118     80'h00_FE00_00_0040_0C8C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2173_1 ( .OUT(na2173_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na2174_2), .IN4(~na532_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2173_2 ( .OUT(na2173_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2173_1_i) );
// C_///AND/      x76y75     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2174_4 ( .OUT(na2174_2), .IN1(1'b1), .IN2(na2173_1), .IN3(na359_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x55y112     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2175_1 ( .OUT(na2175_1_i), .IN1(~na2176_1), .IN2(na536_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2175_2 ( .OUT(na2175_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2175_1_i) );
// C_MX2b////      x49y105     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2176_1 ( .OUT(na2176_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2175_1), .IN7(1'b0), .IN8(~na5888_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x51y121     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2177_1 ( .OUT(na2177_1_i), .IN1(~na2178_1), .IN2(na9255_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2177_2 ( .OUT(na2177_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2177_1_i) );
// C_MX2b////      x55y113     80'h00_0018_00_0040_0A55_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2178_1 ( .OUT(na2178_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_2), .IN4(1'b1), .IN5(~na2177_1), .IN6(1'b0), .IN7(~na5889_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x53y110     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2179_1 ( .OUT(na2179_1_i), .IN1(~na2180_1), .IN2(na9259_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2179_2 ( .OUT(na2179_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2179_1_i) );
// C_MX2b////      x55y69     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2180_1 ( .OUT(na2180_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2179_1), .IN7(1'b0), .IN8(~na5890_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x49y110     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2181_1 ( .OUT(na2181_1_i), .IN1(~na2182_1), .IN2(na9262_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2181_2 ( .OUT(na2181_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2181_1_i) );
// C_MX2b////      x57y81     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2182_1 ( .OUT(na2182_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2181_1), .IN7(1'b0), .IN8(~na5891_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x53y116     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2183_1 ( .OUT(na2183_1_i), .IN1(~na2184_1), .IN2(na9268_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2183_2 ( .OUT(na2183_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2183_1_i) );
// C_MX2b////      x65y85     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2184_1 ( .OUT(na2184_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2183_1), .IN7(1'b0), .IN8(~na5892_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x47y117     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2185_1 ( .OUT(na2185_1_i), .IN1(~na2186_1), .IN2(na582_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2185_2 ( .OUT(na2185_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2185_1_i) );
// C_MX2b////      x59y85     80'h00_0018_00_0040_0A55_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2186_1 ( .OUT(na2186_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_2), .IN4(1'b1), .IN5(~na2185_1), .IN6(1'b0), .IN7(~na5893_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x45y116     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2187_1 ( .OUT(na2187_1_i), .IN1(~na2188_1), .IN2(na9272_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2187_2 ( .OUT(na2187_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2187_1_i) );
// C_MX2b////      x61y89     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2188_1 ( .OUT(na2188_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2187_1), .IN7(1'b0), .IN8(~na5894_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x47y114     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2189_1 ( .OUT(na2189_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2190_1), .IN4(na593_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2189_2 ( .OUT(na2189_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2189_1_i) );
// C_MX2b////      x54y89     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2190_1 ( .OUT(na2190_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2189_1), .IN7(1'b0), .IN8(~na5895_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x51y118     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2191_1 ( .OUT(na2191_1_i), .IN1(~na2192_1), .IN2(na9278_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2191_2 ( .OUT(na2191_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2191_1_i) );
// C_MX2b////      x61y85     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2192_1 ( .OUT(na2192_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2191_1), .IN7(1'b0), .IN8(~na5896_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x50y118     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2193_1 ( .OUT(na2193_1_i), .IN1(~na2194_1), .IN2(na1393_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2193_2 ( .OUT(na2193_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2193_1_i) );
// C_MX2b////      x55y85     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2194_1 ( .OUT(na2194_1), .IN1(1'b1), .IN2(1'b1), .IN3(na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na5897_1), .IN7(1'b0), .IN8(~na2193_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x49y118     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2195_1 ( .OUT(na2195_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2196_1), .IN4(na603_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2195_2 ( .OUT(na2195_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2195_1_i) );
// C_MX2b////      x46y111     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2196_1 ( .OUT(na2196_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2195_1), .IN7(1'b0), .IN8(~na5898_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x49y116     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2197_1 ( .OUT(na2197_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2198_1), .IN4(na609_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2197_2 ( .OUT(na2197_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2197_1_i) );
// C_MX2b////      x50y103     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2198_1 ( .OUT(na2198_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2197_1), .IN7(1'b0), .IN8(~na5899_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x51y120     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2199_1 ( .OUT(na2199_1_i), .IN1(~na2200_1), .IN2(na9287_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2199_2 ( .OUT(na2199_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2199_1_i) );
// C_MX2b////      x47y111     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2200_1 ( .OUT(na2200_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2199_1), .IN7(1'b0), .IN8(~na5900_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x49y112     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2201_1 ( .OUT(na2201_1_i), .IN1(~na2202_1), .IN2(na9284_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2201_2 ( .OUT(na2201_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2201_1_i) );
// C_MX2b////      x47y101     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2202_1 ( .OUT(na2202_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2201_1), .IN7(1'b0), .IN8(~na5901_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x55y114     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2203_1 ( .OUT(na2203_1_i), .IN1(~na2204_1), .IN2(na9290_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2203_2 ( .OUT(na2203_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2203_1_i) );
// C_MX2b////      x49y101     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2204_1 ( .OUT(na2204_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2203_1), .IN7(1'b0), .IN8(~na5902_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x47y110     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2205_1 ( .OUT(na2205_1_i), .IN1(~na2206_1), .IN2(na9524_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2205_2 ( .OUT(na2205_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2205_1_i) );
// C_MX2b////      x45y101     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2206_1 ( .OUT(na2206_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2205_1), .IN7(1'b0), .IN8(~na5903_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x53y114     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2207_1 ( .OUT(na2207_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2208_1), .IN4(na629_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2207_2 ( .OUT(na2207_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2207_1_i) );
// C_MX2b////      x48y103     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2208_1 ( .OUT(na2208_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2207_1), .IN7(1'b0), .IN8(~na5904_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x45y114     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2209_1 ( .OUT(na2209_1_i), .IN1(~na2210_1), .IN2(na9294_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2209_2 ( .OUT(na2209_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2209_1_i) );
// C_MX2b////      x45y107     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2210_1 ( .OUT(na2210_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2209_1), .IN7(1'b0), .IN8(~na5905_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x53y118     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2211_1 ( .OUT(na2211_1_i), .IN1(~na2212_1), .IN2(na9520_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2211_2 ( .OUT(na2211_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2211_1_i) );
// C_MX2b////      x49y107     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2212_1 ( .OUT(na2212_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2211_1), .IN7(1'b0), .IN8(~na5906_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x53y112     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2213_1 ( .OUT(na2213_1_i), .IN1(~na2214_1), .IN2(na9299_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2213_2 ( .OUT(na2213_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2213_1_i) );
// C_MX2b////      x47y103     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2214_1 ( .OUT(na2214_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2213_1), .IN7(1'b0), .IN8(~na5907_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x55y116     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2215_1 ( .OUT(na2215_1_i), .IN1(~na2216_1), .IN2(na9303_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2215_2 ( .OUT(na2215_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2215_1_i) );
// C_MX2b////      x57y111     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2216_1 ( .OUT(na2216_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2215_1), .IN7(1'b0), .IN8(~na5908_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x51y116     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2217_1 ( .OUT(na2217_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2218_1), .IN4(na669_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2217_2 ( .OUT(na2217_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2217_1_i) );
// C_MX2b////      x48y105     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2218_1 ( .OUT(na2218_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2217_1), .IN7(1'b0), .IN8(~na5909_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x55y118     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2219_1 ( .OUT(na2219_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2220_1), .IN4(na674_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2219_2 ( .OUT(na2219_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2219_1_i) );
// C_MX2b////      x52y107     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2220_1 ( .OUT(na2220_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2219_1), .IN7(1'b0), .IN8(~na5910_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x57y114     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2221_1 ( .OUT(na2221_1_i), .IN1(~na2222_1), .IN2(na9307_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2221_2 ( .OUT(na2221_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2221_1_i) );
// C_MX2b////      x51y105     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2222_1 ( .OUT(na2222_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2221_1), .IN7(1'b0), .IN8(~na5911_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x53y120     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2223_1 ( .OUT(na2223_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2224_1), .IN4(na684_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2223_2 ( .OUT(na2223_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2223_1_i) );
// C_MX2b////      x56y117     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2224_1 ( .OUT(na2224_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2223_1), .IN7(1'b0), .IN8(~na5912_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x47y116     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2225_1 ( .OUT(na2225_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2226_1), .IN4(na689_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2225_2 ( .OUT(na2225_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2225_1_i) );
// C_MX2b////      x46y109     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2226_1 ( .OUT(na2226_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2225_1), .IN7(1'b0), .IN8(~na5913_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x53y122     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2227_1 ( .OUT(na2227_1_i), .IN1(~na2228_1), .IN2(na9313_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2227_2 ( .OUT(na2227_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2227_1_i) );
// C_MX2b////      x45y109     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2228_1 ( .OUT(na2228_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2227_1), .IN7(1'b0), .IN8(~na5914_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x57y116     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2229_1 ( .OUT(na2229_1_i), .IN1(~na2230_1), .IN2(na9316_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2229_2 ( .OUT(na2229_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2229_1_i) );
// C_MX2b////      x49y109     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2230_1 ( .OUT(na2230_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2229_1), .IN7(1'b0), .IN8(~na5915_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x55y120     80'h00_FE00_00_0040_0C4C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2231_1 ( .OUT(na2231_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na2232_1), .IN4(na704_1), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2231_2 ( .OUT(na2231_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2231_1_i) );
// C_MX2b////      x58y111     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2232_1 ( .OUT(na2232_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2231_1), .IN7(1'b0), .IN8(~na5916_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x47y118     80'h00_FE00_00_0040_0C13_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2233_1 ( .OUT(na2233_1_i), .IN1(~na2234_1), .IN2(na9321_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3313_2), .IN6(na2172_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2233_2 ( .OUT(na2233_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2233_1_i) );
// C_MX2b////      x47y107     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2234_1 ( .OUT(na2234_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na359_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2233_1), .IN7(1'b0), .IN8(~na5917_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y119     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2235_1 ( .OUT(na2235_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1100_1), .IN6(~na2236_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2235_2 ( .OUT(na2235_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2235_1_i) );
// C_MX2b////      x111y108     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2236_1 ( .OUT(na2236_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1275_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na4005_1), .IN7(1'b0), .IN8(~na1204_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y117     80'h00_FE00_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2237_1 ( .OUT(na2237_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1096_1),
                      .IN8(~na2238_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2237_2 ( .OUT(na2237_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2237_1_i) );
// C_MX2b////      x102y106     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2238_1 ( .OUT(na2238_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1275_1), .IN4(1'b1), .IN5(~na4003_1), .IN6(1'b0), .IN7(~na1202_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x117y95     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2239_1 ( .OUT(na2239_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2239_1), .IN6(na1110_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2239_2 ( .OUT(na2239_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2239_1_i) );
// C_MX4b/D///      x105y117     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2240_1 ( .OUT(na2240_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1094_1), .IN6(~na2241_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2240_2 ( .OUT(na2240_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2240_1_i) );
// C_MX2b////      x111y106     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2241_1 ( .OUT(na2241_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1275_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na4001_2), .IN7(1'b0), .IN8(~na1201_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x108y117     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2242_1 ( .OUT(na2242_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1092_1), .IN6(~na2243_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2242_2 ( .OUT(na2242_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2242_1_i) );
// C_MX2b////      x101y106     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2243_1 ( .OUT(na2243_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1275_1), .IN4(1'b1), .IN5(~na3998_2), .IN6(1'b0), .IN7(~na9447_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x106y120     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2244_1 ( .OUT(na2244_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1090_1), .IN6(~na2245_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2244_2 ( .OUT(na2244_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2244_1_i) );
// C_MX2b////      x111y90     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2245_1 ( .OUT(na2245_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1275_1), .IN4(1'b1), .IN5(~na3998_1), .IN6(1'b0), .IN7(~na9445_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x119y85     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2246_1 ( .OUT(na2246_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1095_2),
                      .IN8(na9567_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2246_2 ( .OUT(na2246_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2246_1_i) );
// C_AND////      x122y65     80'h00_0018_00_0000_0C88_42FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2248_1 ( .OUT(na2248_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3290_1), .IN6(~na9801_2), .IN7(~na3596_2),
                      .IN8(na983_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x129y54     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2249_1 ( .OUT(na2249_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na500_2), .IN5(1'b0), .IN6(~na2718_2), .IN7(1'b0), .IN8(~na7889_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x130y53     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2250_1 ( .OUT(na2250_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2746_2), .IN6(na2718_1), .IN7(na2737_1),
                      .IN8(na9665_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x105y110     80'h00_FE00_00_0040_0A3C_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2251_1 ( .OUT(na2251_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na2251_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2251_2 ( .OUT(na2251_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2251_1_i) );
// C_AND/D///      x87y74     80'h00_FE00_00_0000_0888_F128
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2252_1 ( .OUT(na2252_1_i), .IN1(na468_1), .IN2(na27_1), .IN3(na469_1), .IN4(~na6626_1), .IN5(~na32_1), .IN6(~na2252_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2252_2 ( .OUT(na2252_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2252_1_i) );
// C_MX4b/D///      x107y99     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2253_1 ( .OUT(na2253_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2253_1), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2253_2 ( .OUT(na2253_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2253_1_i) );
// C_MX4b/D///      x123y85     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2254_1 ( .OUT(na2254_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2254_1), .IN6(na993_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2254_2 ( .OUT(na2254_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2254_1_i) );
// C_MX4b/D///      x98y108     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2255_1 ( .OUT(na2255_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3764_1),
                      .IN8(na2255_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2255_2 ( .OUT(na2255_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2255_1_i) );
// C_MX2b/D///      x67y117     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2256_1 ( .OUT(na2256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na404_1), .IN5(1'b0), .IN6(na46_1), .IN7(1'b0), .IN8(na520_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2256_2 ( .OUT(na2256_1), .CLK(na4116_1), .EN(~na359_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2256_1_i) );
// C_AND////      x68y51     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2257_1 ( .OUT(na2257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b1), .IN8(na5961_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x59y68     80'h00_0018_00_0000_0CEE_5C00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2262_1 ( .OUT(na2262_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na7890_2), .IN7(~na2263_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y63     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2263_1 ( .OUT(na2263_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na9802_2), .IN5(1'b0), .IN6(~na5948_1), .IN7(1'b0), .IN8(~na7891_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x58y89     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2264_1 ( .OUT(na2264_1), .IN1(na5972_1), .IN2(na5953_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x56y66     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2265_1 ( .OUT(na2265_1), .IN1(na5972_1), .IN2(na5953_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x57y65     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2266_1 ( .OUT(na2266_1), .IN1(na5972_1), .IN2(na9913_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x63y65     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2267_1 ( .OUT(na2267_1), .IN1(na5972_1), .IN2(na5956_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x61y66     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2268_1 ( .OUT(na2268_1), .IN1(na5972_1), .IN2(na5957_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x65y67     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2269_1 ( .OUT(na2269_1), .IN1(na5972_1), .IN2(na9914_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x65y66     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2270_1 ( .OUT(na2270_1), .IN1(na5972_1), .IN2(na5959_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x68y70     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2271_1 ( .OUT(na2271_1), .IN1(na5972_1), .IN2(na5960_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x57y64     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2272_4 ( .OUT(na2272_2), .IN1(na3329_2), .IN2(na3263_1), .IN3(na5263_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x62y57     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2273_4 ( .OUT(na2273_2), .IN1(na3329_2), .IN2(na3263_1), .IN3(na5264_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x56y63     80'h00_0018_00_0040_0C0C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2274_1 ( .OUT(na2274_1), .IN1(1'b0), .IN2(1'b0), .IN3(na6308_1), .IN4(na5265_1), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x56y59     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2275_1 ( .OUT(na2275_1), .IN1(na9938_2), .IN2(na5266_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x68y64     80'h00_0018_00_0040_0C0C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2276_1 ( .OUT(na2276_1), .IN1(1'b0), .IN2(1'b0), .IN3(na9939_2), .IN4(na5267_1), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x74y74     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2277_1 ( .OUT(na2277_1), .IN1(na6324_2), .IN2(na5268_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x68y65     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2278_1 ( .OUT(na2278_1), .IN1(na6312_2), .IN2(na5269_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x61y67     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2279_1 ( .OUT(na2279_1), .IN1(na6313_1), .IN2(na5270_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x57y66     80'h00_0018_00_0040_0C0C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2280_1 ( .OUT(na2280_1), .IN1(1'b0), .IN2(1'b0), .IN3(na6314_2), .IN4(na5271_1), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y65     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2281_1 ( .OUT(na2281_1), .IN1(na6315_1), .IN2(na5272_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x56y58     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2282_1 ( .OUT(na2282_1), .IN1(na6325_2), .IN2(na5273_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x70y53     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2283_1 ( .OUT(na2283_1), .IN1(na6317_2), .IN2(na5274_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x59y62     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2284_1 ( .OUT(na2284_1), .IN1(na6318_1), .IN2(na5275_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x53y72     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2285_1 ( .OUT(na2285_1), .IN1(na6319_2), .IN2(na5276_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y59     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2286_1 ( .OUT(na2286_1), .IN1(na6320_1), .IN2(na5277_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y61     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2287_1 ( .OUT(na2287_1), .IN1(na6321_1), .IN2(na5278_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y64     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2288_1 ( .OUT(na2288_1), .IN1(na6322_2), .IN2(na5279_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y67     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2289_1 ( .OUT(na2289_1), .IN1(na6323_1), .IN2(na5280_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x56y70     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2290_1 ( .OUT(na2290_1), .IN1(na6324_1), .IN2(na5281_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x55y68     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2291_1 ( .OUT(na2291_1), .IN1(na6325_1), .IN2(na5282_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y69     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2292_1 ( .OUT(na2292_1), .IN1(na6326_2), .IN2(na5283_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y75     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2293_1 ( .OUT(na2293_1), .IN1(na6327_1), .IN2(na5284_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y73     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2294_1 ( .OUT(na2294_1), .IN1(na6328_2), .IN2(na5285_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x50y71     80'h00_0018_00_0040_0C0C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2295_1 ( .OUT(na2295_1), .IN1(1'b0), .IN2(1'b0), .IN3(na6329_1), .IN4(na5286_1), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y74     80'h00_0018_00_0040_0C0C_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2296_1 ( .OUT(na2296_1), .IN1(1'b0), .IN2(1'b0), .IN3(na6330_2), .IN4(na5287_1), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x56y55     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2297_1 ( .OUT(na2297_1), .IN1(na6331_1), .IN2(na5288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y62     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2298_1 ( .OUT(na2298_1), .IN1(na6332_2), .IN2(na5289_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x48y55     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2299_1 ( .OUT(na2299_1), .IN1(na6333_1), .IN2(na5290_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y58     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2300_1 ( .OUT(na2300_1), .IN1(na6334_2), .IN2(na5291_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x52y78     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2301_1 ( .OUT(na2301_1), .IN1(na6335_1), .IN2(na5292_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x64y79     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2302_1 ( .OUT(na2302_1), .IN1(na6336_2), .IN2(na5293_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x50y59     80'h00_0018_00_0040_0C03_0800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2303_1 ( .OUT(na2303_1), .IN1(na6320_2), .IN2(na5294_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(na3263_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y79     80'h00_0018_00_0000_0888_4C14
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2306_1 ( .OUT(na2306_1), .IN1(~na9574_2), .IN2(na7893_1), .IN3(~na2321_1), .IN4(~na2322_1), .IN5(1'b1), .IN6(na9573_2), .IN7(~na2318_1),
                      .IN8(na2322_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x59y71     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2309_1 ( .OUT(na2309_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2310_1), .IN6(na7895_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2309_4 ( .OUT(na2309_2), .IN1(na554_2), .IN2(na5270_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x67y65     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2310_1 ( .OUT(na2310_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5256_1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x56y68     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2311_1 ( .OUT(na2311_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7897_1), .IN7(1'b1), .IN8(na2312_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x70y70     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2312_1 ( .OUT(na2312_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5255_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y70     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2314_4 ( .OUT(na2314_2), .IN1(1'b1), .IN2(na2315_1), .IN3(na7899_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x67y70     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2315_1 ( .OUT(na2315_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na9879_2), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y69     80'h00_0078_00_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2316_1 ( .OUT(na2316_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7901_1), .IN7(1'b1), .IN8(na2317_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2316_4 ( .OUT(na2316_2), .IN1(na554_2), .IN2(na5274_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y42     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2317_1 ( .OUT(na2317_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na5250_1), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x54y79     80'h00_0078_00_0000_0C66_5A60
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2318_1 ( .OUT(na2318_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2378_2), .IN6(1'b0), .IN7(~na2316_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2318_4 ( .OUT(na2318_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2316_1), .IN4(na667_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x54y81     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2320_1 ( .OUT(na2320_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na9872_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x62y81     80'h00_0078_00_0000_0C66_5AA3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2321_1 ( .OUT(na2321_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na540_1), .IN6(1'b0), .IN7(~na3491_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2321_4 ( .OUT(na2321_2), .IN1(1'b0), .IN2(~na2314_2), .IN3(na661_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x50y68     80'h00_0078_00_0000_0C66_A5AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2322_1 ( .OUT(na2322_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2309_2), .IN6(1'b0), .IN7(na589_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2322_4 ( .OUT(na2322_2), .IN1(na2309_1), .IN2(1'b0), .IN3(na9315_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x74y69     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2324_1 ( .OUT(na2324_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na9928_2), .IN6(~na5235_1), .IN7(1'b1),
                      .IN8(~na5969_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x51y70     80'h00_0018_00_0000_0888_6666
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2325_1 ( .OUT(na2325_1), .IN1(na687_1), .IN2(~na9576_2), .IN3(na637_1), .IN4(~na9578_2), .IN5(na9256_2), .IN6(~na3489_1),
                      .IN7(~na2327_2), .IN8(na9579_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x52y71     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2327_1 ( .OUT(na2327_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2328_1), .IN6(na7910_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2327_4 ( .OUT(na2327_2), .IN1(na554_2), .IN2(na5273_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y45     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2328_1 ( .OUT(na2328_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5254_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y58     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2331_1 ( .OUT(na2331_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5971_1), .IN6(1'b1), .IN7(~na5238_2),
                      .IN8(~na9931_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x57y67     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2332_1 ( .OUT(na2332_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7912_2), .IN6(na2333_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2332_4 ( .OUT(na2332_2), .IN1(na7912_1), .IN2(na2331_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y42     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2333_1 ( .OUT(na2333_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na5247_2), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x61y65     80'h00_0018_00_0000_0C88_66FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2334_1 ( .OUT(na2334_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3487_1), .IN6(na9261_2), .IN7(na2335_2),
                      .IN8(~na594_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x68y63     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2335_4 ( .OUT(na2335_2), .IN1(na7918_2), .IN2(1'b1), .IN3(na2336_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y65     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2336_1 ( .OUT(na2336_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5971_2), .IN6(1'b1), .IN7(~na5237_1),
                      .IN8(~na9932_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x66y62     80'h00_0060_00_0000_0C08_FF66
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2337_4 ( .OUT(na2337_2), .IN1(na2338_2), .IN2(~na9274_2), .IN3(~na9583_2), .IN4(na682_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y65     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2338_4 ( .OUT(na2338_2), .IN1(1'b1), .IN2(na2339_1), .IN3(na7922_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y60     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2339_1 ( .OUT(na2339_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na9926_2), .IN6(1'b1), .IN7(~na9867_2),
                      .IN8(~na5969_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x55y70     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2340_4 ( .OUT(na2340_2), .IN1(na2341_1), .IN2(1'b1), .IN3(na7924_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y39     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2341_1 ( .OUT(na2341_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na9883_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x53y69     80'h00_0018_00_0000_0888_4141
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2342_1 ( .OUT(na2342_1), .IN1(~na2361_1), .IN2(~na2364_1), .IN3(~na2344_1), .IN4(na7934_1), .IN5(~na2361_2), .IN6(~na2364_2),
                      .IN7(~na2344_2), .IN8(na7934_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x56y77     80'h00_0078_00_0000_0C66_A5C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2344_1 ( .OUT(na2344_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2354_2), .IN6(1'b0), .IN7(na723_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2344_4 ( .OUT(na2344_2), .IN1(~na2354_1), .IN2(1'b0), .IN3(1'b0), .IN4(na622_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y39     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2346_1 ( .OUT(na2346_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na9889_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y64     80'h00_0078_00_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2348_1 ( .OUT(na2348_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7928_1), .IN6(na2349_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2348_4 ( .OUT(na2348_2), .IN1(na554_2), .IN2(na5269_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y42     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2349_1 ( .OUT(na2349_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5252_1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x57y69     80'h00_0078_00_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2351_1 ( .OUT(na2351_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7930_2), .IN6(1'b1), .IN7(na2352_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2351_4 ( .OUT(na2351_2), .IN1(na2366_1), .IN2(na7942_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y39     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2352_1 ( .OUT(na2352_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na5258_1), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x51y69     80'h00_0078_00_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2354_1 ( .OUT(na2354_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7926_2), .IN6(na2355_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2354_4 ( .OUT(na2354_2), .IN1(na7926_1), .IN2(1'b1), .IN3(na2346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y46     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2355_1 ( .OUT(na2355_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na9875_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y75     80'h00_0078_00_0000_0C88_CACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2357_1 ( .OUT(na2357_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7936_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2358_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2357_4 ( .OUT(na2357_2), .IN1(1'b1), .IN2(na7938_2), .IN3(1'b1), .IN4(na2360_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y38     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2358_1 ( .OUT(na2358_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na5248_1), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y44     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2360_1 ( .OUT(na2360_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5241_1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y71     80'h00_0078_00_0000_0C66_3A90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2361_1 ( .OUT(na2361_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2362_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na2348_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2361_4 ( .OUT(na2361_2), .IN1(1'b0), .IN2(1'b0), .IN3(na677_1), .IN4(~na2348_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x57y63     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2362_1 ( .OUT(na2362_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7940_2), .IN6(1'b1), .IN7(na2363_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y53     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2363_1 ( .OUT(na2363_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5967_1), .IN6(1'b1), .IN7(~na5234_2),
                      .IN8(~na9924_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x57y78     80'h00_0078_00_0000_0C66_A5A5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2364_1 ( .OUT(na2364_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2351_2), .IN6(1'b0), .IN7(na672_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2364_4 ( .OUT(na2364_2), .IN1(~na2351_1), .IN2(1'b0), .IN3(na707_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y37     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2366_1 ( .OUT(na2366_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na9881_2), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x47y60     80'h00_0018_00_0000_0888_6666
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2367_1 ( .OUT(na2367_1), .IN1(na1603_1), .IN2(~na9588_2), .IN3(na632_1), .IN4(~na2372_1), .IN5(~na2378_1), .IN6(na9281_2),
                      .IN7(~na2369_2), .IN8(na2372_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y73     80'h00_0078_00_0000_0C88_8FF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2369_1 ( .OUT(na2369_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2370_1), .IN8(na7944_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2369_4 ( .OUT(na2369_2), .IN1(na554_2), .IN2(na5268_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y43     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2370_1 ( .OUT(na2370_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5245_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y76     80'h00_0078_00_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2372_1 ( .OUT(na2372_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2373_1), .IN7(na7948_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2372_4 ( .OUT(na2372_2), .IN1(1'b1), .IN2(na2376_1), .IN3(na7948_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y44     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2373_1 ( .OUT(na2373_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5246_1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y52     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2376_1 ( .OUT(na2376_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5967_2), .IN6(~na5233_1), .IN7(1'b1),
                      .IN8(~na9925_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x47y55     80'h00_0078_00_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2378_1 ( .OUT(na2378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2379_1), .IN7(1'b1), .IN8(na7950_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2378_4 ( .OUT(na2378_2), .IN1(1'b1), .IN2(na7903_1), .IN3(na2320_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y44     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2379_1 ( .OUT(na2379_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na9873_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y55     80'h00_0018_00_0000_0888_F88C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2380_1 ( .OUT(na2380_1), .IN1(1'b1), .IN2(na7953_2), .IN3(na7952_2), .IN4(na7954_1), .IN5(na7955_1), .IN6(na7953_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x53y79     80'h00_0078_00_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2383_1 ( .OUT(na2383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2384_1), .IN7(1'b1), .IN8(na7957_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2383_4 ( .OUT(na2383_2), .IN1(1'b1), .IN2(na7961_1), .IN3(1'b1), .IN4(na2388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y40     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2384_1 ( .OUT(na2384_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na5244_1), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y81     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2385_1 ( .OUT(na2385_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7959_1), .IN7(na2386_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y41     80'h00_0018_00_0040_0ADF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2386_1 ( .OUT(na2386_1), .IN1(1'b1), .IN2(na369_2), .IN3(~na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(1'b1), .IN7(~na5257_2),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y42     80'h00_0018_00_0040_0ABF_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2388_1 ( .OUT(na2388_1), .IN1(1'b1), .IN2(~na369_2), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5972_1), .IN6(~na9877_2), .IN7(1'b1),
                      .IN8(~na9933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y77     80'h00_0018_00_0040_0AF7_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2389_1 ( .OUT(na2389_1), .IN1(na2354_2), .IN2(1'b1), .IN3(na723_1), .IN4(1'b1), .IN5(~na3269_2), .IN6(~na9594_2), .IN7(~na2390_1),
                      .IN8(na9807_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x64y77     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2390_1 ( .OUT(na2390_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na723_1), .IN8(na6367_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2390_5 ( .OUT(na2390_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2390_1) );
// C_MX2b////      x55y79     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2391_1 ( .OUT(na2391_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2596_1), .IN8(na355_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y83     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2392_1 ( .OUT(na2392_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1377_1), .IN5(na540_1), .IN6(1'b0), .IN7(na2597_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y90     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2393_1 ( .OUT(na2393_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na9633_2), .IN6(1'b0), .IN7(na545_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x57y88     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2394_1 ( .OUT(na2394_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na2599_1), .IN6(1'b0), .IN7(na550_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x58y81     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2395_1 ( .OUT(na2395_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2369_2), .IN8(na9634_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x57y79     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2396_1 ( .OUT(na2396_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2601_1), .IN8(na2348_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y88     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2397_1 ( .OUT(na2397_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2309_2), .IN6(na9636_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y85     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2398_1 ( .OUT(na2398_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na589_1), .IN8(na9637_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y87     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2399_1 ( .OUT(na2399_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2604_1), .IN8(na594_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y89     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2400_1 ( .OUT(na2400_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na2605_1), .IN6(1'b0), .IN7(na2327_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y86     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2401_1 ( .OUT(na2401_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na2606_1), .IN6(1'b0), .IN7(na2316_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y96     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2402_1 ( .OUT(na2402_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na607_1), .IN8(na2607_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y93     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2403_1 ( .OUT(na2403_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1377_1), .IN5(1'b0), .IN6(na2608_1), .IN7(1'b0), .IN8(na612_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y91     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2404_1 ( .OUT(na2404_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9639_2), .IN8(na622_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y90     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2405_1 ( .OUT(na2405_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2610_1), .IN8(na617_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y88     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2406_1 ( .OUT(na2406_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na627_1), .IN8(na2611_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y89     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2407_1 ( .OUT(na2407_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1377_1), .IN5(na1603_1), .IN6(1'b0), .IN7(na2612_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y91     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2408_1 ( .OUT(na2408_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na9641_2), .IN6(1'b0), .IN7(na632_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x51y93     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2409_1 ( .OUT(na2409_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na637_1), .IN8(na2614_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x57y94     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2410_1 ( .OUT(na2410_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1586_1), .IN6(na9642_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y94     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2411_1 ( .OUT(na2411_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na9643_2), .IN6(1'b0), .IN7(na661_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x59y95     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2412_1 ( .OUT(na2412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1377_1), .IN5(1'b0), .IN6(na2617_1), .IN7(1'b0), .IN8(na667_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y93     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2413_1 ( .OUT(na2413_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na2618_1), .IN6(1'b0), .IN7(na672_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x51y96     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2414_1 ( .OUT(na2414_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na2619_1), .IN6(1'b0), .IN7(na677_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y94     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2415_1 ( .OUT(na2415_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2620_1), .IN8(na682_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y95     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2416_1 ( .OUT(na2416_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b0), .IN4(1'b0), .IN5(na687_1), .IN6(na2621_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y95     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2417_1 ( .OUT(na2417_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na2622_1), .IN6(1'b0), .IN7(na692_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x57y96     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2418_1 ( .OUT(na2418_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1377_1), .IN5(na697_1), .IN6(1'b0), .IN7(na2623_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y95     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2419_1 ( .OUT(na2419_1), .IN1(1'b1), .IN2(~na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2624_1), .IN8(na702_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x57y95     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2420_1 ( .OUT(na2420_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1377_1), .IN5(na2625_1), .IN6(1'b0), .IN7(na707_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x58y94     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2421_1 ( .OUT(na2421_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na723_1), .IN8(na9647_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b*////D      x52y80     80'h00_FA18_00_0040_0531_000C
C_MX2b     #(.CPE_CFG (9'b1_0000_0000)) 
           _a2422_1 ( .OUT(na2422_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na50_1), .IN6(na9603_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2422_5 ( .OUT(na2422_2), .CLK(na4116_1), .EN(na347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2422_1) );
// C_MX2b////D      x62y65     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2423_1 ( .OUT(na2423_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na540_1), .IN6(1'b0), .IN7(na6354_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2423_5 ( .OUT(na2423_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2423_1) );
// C_MX2b////D      x66y71     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2424_1 ( .OUT(na2424_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na545_1), .IN8(na6368_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2424_5 ( .OUT(na2424_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2424_1) );
// C_MX2b////D      x52y68     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2425_1 ( .OUT(na2425_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na550_1), .IN8(na6368_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2425_5 ( .OUT(na2425_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2425_1) );
// C_MX2b////D      x62y68     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2426_1 ( .OUT(na2426_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na9589_2), .IN6(1'b0), .IN7(na6370_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2426_5 ( .OUT(na2426_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2426_1) );
// C_MX2b////D      x55y65     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2427_1 ( .OUT(na2427_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6370_2), .IN8(na2348_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2427_5 ( .OUT(na2427_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2427_1) );
// C_MX2b////D      x56y65     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2428_1 ( .OUT(na2428_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9568_2), .IN8(na6372_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2428_5 ( .OUT(na2428_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2428_1) );
// C_MX2b////D      x59y70     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2429_1 ( .OUT(na2429_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na589_1), .IN8(na6372_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2429_5 ( .OUT(na2429_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2429_1) );
// C_MX2b////D      x53y71     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2430_1 ( .OUT(na2430_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6374_1), .IN8(na594_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2430_5 ( .OUT(na2430_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2430_1) );
// C_MX2b////D      x61y73     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2431_1 ( .OUT(na2431_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na9577_2), .IN6(1'b0), .IN7(na6374_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2431_5 ( .OUT(na2431_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2431_1) );
// C_MX2b////D      x55y67     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2432_1 ( .OUT(na2432_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2316_2), .IN8(na6345_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2432_5 ( .OUT(na2432_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2432_1) );
// C_MX2b////D      x61y74     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2433_1 ( .OUT(na2433_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na607_1), .IN8(na6345_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2433_5 ( .OUT(na2433_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2433_1) );
// C_MX2b////D      x63y72     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2434_1 ( .OUT(na2434_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6347_1), .IN8(na612_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2434_5 ( .OUT(na2434_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2434_1) );
// C_MX2b////D      x63y73     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2435_1 ( .OUT(na2435_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6347_2), .IN8(na622_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2435_5 ( .OUT(na2435_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2435_1) );
// C_MX2b////D      x63y67     80'h00_F618_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2436_1 ( .OUT(na2436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na9821_2), .IN5(1'b0), .IN6(na9286_2), .IN7(1'b0), .IN8(na6349_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2436_5 ( .OUT(na2436_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2436_1) );
// C_MX2b////D      x73y74     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2437_1 ( .OUT(na2437_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na627_1), .IN8(na6349_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2437_5 ( .OUT(na2437_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2437_1) );
// C_MX2b////D      x71y76     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2438_1 ( .OUT(na2438_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na1603_1), .IN6(1'b0), .IN7(na6351_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2438_5 ( .OUT(na2438_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2438_1) );
// C_MX2b////D      x72y76     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2439_1 ( .OUT(na2439_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na9292_2), .IN6(1'b0), .IN7(na6351_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2439_5 ( .OUT(na2439_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2439_1) );
// C_MX2b////D      x71y75     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2440_1 ( .OUT(na2440_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na637_1), .IN8(na6353_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2440_5 ( .OUT(na2440_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2440_1) );
// C_MX2b////D      x70y79     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2441_1 ( .OUT(na2441_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9522_2), .IN8(na6353_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2441_5 ( .OUT(na2441_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2441_1) );
// C_MX2b////D      x86y79     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2442_1 ( .OUT(na2442_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na9301_2), .IN6(1'b0), .IN7(na6356_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2442_5 ( .OUT(na2442_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2442_1) );
// C_MX2b////D      x88y61     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2443_1 ( .OUT(na2443_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6356_2), .IN8(na667_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2443_5 ( .OUT(na2443_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2443_1) );
// C_MX2b////D      x66y75     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2444_1 ( .OUT(na2444_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na672_1), .IN8(na6358_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2444_5 ( .OUT(na2444_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2444_1) );
// C_MX2b////D      x70y69     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2445_1 ( .OUT(na2445_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na677_1), .IN8(na6358_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2445_5 ( .OUT(na2445_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2445_1) );
// C_MX2b////D      x60y76     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2446_1 ( .OUT(na2446_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6360_1), .IN8(na682_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2446_5 ( .OUT(na2446_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2446_1) );
// C_MX2b////D      x66y86     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2447_1 ( .OUT(na2447_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na687_1), .IN6(1'b0), .IN7(na6360_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2447_5 ( .OUT(na2447_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2447_1) );
// C_MX2b////D      x62y79     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2448_1 ( .OUT(na2448_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na692_1), .IN8(na6362_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2448_5 ( .OUT(na2448_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2448_1) );
// C_MX2b////D      x68y77     80'h00_F618_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2449_1 ( .OUT(na2449_1), .IN1(1'b1), .IN2(~na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9315_2), .IN8(na6362_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2449_5 ( .OUT(na2449_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2449_1) );
// C_MX2b////D      x66y78     80'h00_F618_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2450_1 ( .OUT(na2450_1), .IN1(1'b1), .IN2(na3330_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6364_1), .IN8(na702_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2450_5 ( .OUT(na2450_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2450_1) );
// C_MX2b////D      x67y77     80'h00_F618_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2451_1 ( .OUT(na2451_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9821_2), .IN5(na9318_2), .IN6(1'b0), .IN7(na6364_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2451_5 ( .OUT(na2451_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2451_1) );
// C_MX4b////      x65y58     80'h00_0018_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2454_1 ( .OUT(na2454_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na9908_2), .IN6(~na3585_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y61     80'h00_0018_00_0040_0A31_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2455_1 ( .OUT(na2455_1), .IN1(~na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(~na2456_1), .IN6(na5706_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x65y59     80'h00_0078_00_0000_0C88_53CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2456_1 ( .OUT(na2456_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2457_2), .IN7(~na7963_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2456_4 ( .OUT(na2456_2), .IN1(na1372_1), .IN2(1'b1), .IN3(1'b1), .IN4(na5974_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y58     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2457_4 ( .OUT(na2457_2), .IN1(~na5692_2), .IN2(~na3585_1), .IN3(~na5925_2), .IN4(~na9906_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y60     80'h00_0018_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2459_1 ( .OUT(na2459_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na5705_2), .IN5(1'b0), .IN6(1'b0), .IN7(na5707_2),
                      .IN8(~na2460_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x76y58     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2460_4 ( .OUT(na2460_2), .IN1(~na7967_1), .IN2(~na2457_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y58     80'h00_0018_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2462_1 ( .OUT(na2462_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5708_2), .IN6(~na2463_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x71y60     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2463_4 ( .OUT(na2463_2), .IN1(1'b1), .IN2(~na2457_2), .IN3(1'b1), .IN4(~na7971_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y60     80'h00_0018_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2465_1 ( .OUT(na2465_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5709_2), .IN6(~na2466_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x75y62     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2466_1 ( .OUT(na2466_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9613_2), .IN6(~na7975_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y61     80'h00_0018_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2468_1 ( .OUT(na2468_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na5705_2), .IN5(1'b0), .IN6(1'b0), .IN7(na5710_1),
                      .IN8(~na2469_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y56     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2469_4 ( .OUT(na2469_2), .IN1(1'b1), .IN2(~na2457_2), .IN3(1'b1), .IN4(~na7979_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y67     80'h00_0018_00_0040_0A31_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2471_1 ( .OUT(na2471_1), .IN1(~na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(~na2472_2), .IN6(na5711_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y63     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2472_4 ( .OUT(na2472_2), .IN1(1'b1), .IN2(~na2457_2), .IN3(1'b1), .IN4(~na7983_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x62y59     80'h00_0018_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2474_1 ( .OUT(na2474_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na5705_2), .IN5(1'b0), .IN6(1'b0), .IN7(na5712_2),
                      .IN8(~na2475_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y58     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2475_1 ( .OUT(na2475_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2457_2), .IN7(1'b1), .IN8(~na7987_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x70y68     80'h00_0018_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2477_1 ( .OUT(na2477_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5713_1), .IN6(~na2478_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x73y60     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2478_1 ( .OUT(na2478_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na2457_2), .IN7(na10016_2), .IN8(na2479_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y62     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2479_1 ( .OUT(na2479_1), .IN1(na7966_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9552_2), .IN8(~na2148_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x73y68     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2480_1 ( .OUT(na2480_1), .IN1(na7994_2), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5714_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y64     80'h00_0060_00_0000_0C08_FF52
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2481_4 ( .OUT(na2481_2), .IN1(na2456_2), .IN2(~na2457_2), .IN3(~na2482_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y69     80'h00_0018_00_0000_0C88_14FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2482_1 ( .OUT(na2482_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na5692_2), .IN6(na9905_2), .IN7(~na5925_2),
                      .IN8(~na2479_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x62y61     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2484_1 ( .OUT(na2484_1), .IN1(na7997_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5715_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x68y42     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2486_1 ( .OUT(na2486_1), .IN1(na8000_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5716_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x67y45     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2488_1 ( .OUT(na2488_1), .IN1(na8003_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5717_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x72y57     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2490_1 ( .OUT(na2490_1), .IN1(na8006_2), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5718_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x70y57     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2492_1 ( .OUT(na2492_1), .IN1(na8009_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5719_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x67y57     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2494_1 ( .OUT(na2494_1), .IN1(na8012_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5720_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x65y57     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2496_1 ( .OUT(na2496_1), .IN1(na8015_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5721_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x74y57     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2498_1 ( .OUT(na2498_1), .IN1(na8018_2), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5722_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x74y56     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2500_1 ( .OUT(na2500_1), .IN1(na8021_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5723_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x72y44     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2502_1 ( .OUT(na2502_1), .IN1(na8024_2), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5724_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x69y39     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2504_1 ( .OUT(na2504_1), .IN1(na8027_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5725_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x72y46     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2506_1 ( .OUT(na2506_1), .IN1(na8030_2), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5726_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x71y47     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2508_1 ( .OUT(na2508_1), .IN1(na8033_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5727_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x72y48     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2510_1 ( .OUT(na2510_1), .IN1(na8036_2), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5728_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x70y40     80'h00_0018_00_0000_0888_FE3B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2512_1 ( .OUT(na2512_1), .IN1(na8039_1), .IN2(~na2481_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(na2456_2), .IN6(na5729_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y59     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2514_4 ( .OUT(na2514_2), .IN1(1'b1), .IN2(1'b1), .IN3(na5684_2), .IN4(~na5705_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y58     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2515_4 ( .OUT(na2515_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na9909_2), .IN4(na5685_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x62y62     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2516_1 ( .OUT(na2516_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5686_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na5705_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x61y61     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2517_1 ( .OUT(na2517_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5687_2), .IN7(1'b1), .IN8(~na5705_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x56y56     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2518_4 ( .OUT(na2518_2), .IN1(1'b1), .IN2(1'b1), .IN3(na5688_2), .IN4(~na5705_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x68y66     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2519_4 ( .OUT(na2519_2), .IN1(~na1372_1), .IN2(~na9502_2), .IN3(1'b0), .IN4(~na5705_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x67y75     80'h00_F600_80_0000_0C07_FFA7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a2520_4 ( .OUT(na2520_2_i), .IN1(~na5236_2), .IN2(~na5953_2), .IN3(na2521_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2520_5 ( .OUT(na2520_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2520_2_i) );
// C_MX4b////      x74y67     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2521_1 ( .OUT(na2521_1), .IN1(1'b1), .IN2(na5953_1), .IN3(1'b1), .IN4(~na9912_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na5228_2),
                      .IN8(~na9868_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x67y75     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2522_1 ( .OUT(na2522_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9869_2), .IN6(~na5953_2), .IN7(na2523_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2522_2 ( .OUT(na2522_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2522_1_i) );
// C_MX4b////      x72y81     80'h00_0018_00_0040_0A3F_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2523_1 ( .OUT(na2523_1), .IN1(1'b1), .IN2(na5953_1), .IN3(1'b1), .IN4(na9912_2), .IN5(~na5229_1), .IN6(~na9870_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x69y78     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2524_1 ( .OUT(na2524_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9871_2), .IN6(~na5953_2), .IN7(na2525_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2524_2 ( .OUT(na2524_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2524_1_i) );
// C_MX4b////      x72y79     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2525_1 ( .OUT(na2525_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b1), .IN4(~na9912_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na5238_2),
                      .IN8(~na5230_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x68y68     80'h00_F600_80_0000_0C07_FFC7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a2526_4 ( .OUT(na2526_2_i), .IN1(~na5239_2), .IN2(~na5953_2), .IN3(1'b0), .IN4(na2527_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2526_5 ( .OUT(na2526_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2526_2_i) );
// C_MX4b////      x68y78     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2527_1 ( .OUT(na2527_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b1), .IN4(~na9912_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na9872_2),
                      .IN8(~na5231_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x70y72     80'h00_F600_80_0000_0C07_FFC7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a2528_4 ( .OUT(na2528_2_i), .IN1(~na5240_1), .IN2(~na5953_2), .IN3(1'b0), .IN4(na2529_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2528_5 ( .OUT(na2528_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2528_2_i) );
// C_MX4b////      x76y76     80'h00_0018_00_0040_0ACF_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2529_1 ( .OUT(na2529_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b1), .IN4(~na9912_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na9873_2),
                      .IN8(~na5232_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x72y70     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2530_1 ( .OUT(na2530_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9874_2), .IN6(~na5953_2), .IN7(na2531_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2530_2 ( .OUT(na2530_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2530_1_i) );
// C_MX4b////      x72y75     80'h00_0018_00_0040_0A3F_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2531_1 ( .OUT(na2531_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b1), .IN4(na9912_2), .IN5(~na9874_2), .IN6(~na5233_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x74y72     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2532_1 ( .OUT(na2532_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na5242_1), .IN6(~na5953_2), .IN7(na2533_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2532_2 ( .OUT(na2532_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2532_1_i) );
// C_MX4b////      x74y79     80'h00_0018_00_0040_0ACF_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2533_1 ( .OUT(na2533_1), .IN1(1'b1), .IN2(na5953_1), .IN3(1'b1), .IN4(~na9912_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na5234_2),
                      .IN8(~na9876_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x78y73     80'h00_F600_80_0000_0C07_FFA7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a2534_4 ( .OUT(na2534_2_i), .IN1(~na5243_2), .IN2(~na5953_2), .IN3(na2535_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2534_5 ( .OUT(na2534_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2534_2_i) );
// C_MX4b////      x80y73     80'h00_0018_00_0040_0A3F_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2535_1 ( .OUT(na2535_1), .IN1(1'b1), .IN2(~na5953_1), .IN3(1'b1), .IN4(na9912_2), .IN5(~na5243_2), .IN6(~na5235_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x76y70     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2536_1 ( .OUT(na2536_1_i), .IN1(1'b1), .IN2(na5953_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na5228_2), .IN8(na9878_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2536_2 ( .OUT(na2536_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2536_1_i) );
// C_MX2b/D///      x71y71     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2537_1 ( .OUT(na2537_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na9912_2), .IN5(na5229_1), .IN6(1'b0), .IN7(na5245_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2537_2 ( .OUT(na2537_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2537_1_i) );
// C_MX2b/D///      x72y63     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2538_1 ( .OUT(na2538_1_i), .IN1(1'b1), .IN2(~na5953_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na5246_1), .IN8(na5230_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2538_2 ( .OUT(na2538_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2538_1_i) );
// C_MX2b/D///      x72y65     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2539_1 ( .OUT(na2539_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na9912_2), .IN5(1'b0), .IN6(na5247_2), .IN7(1'b0), .IN8(na5231_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2539_2 ( .OUT(na2539_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2539_1_i) );
// C_MX2b/D///      x71y63     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2540_1 ( .OUT(na2540_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na9912_2), .IN5(1'b0), .IN6(na5248_1), .IN7(1'b0), .IN8(na5232_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2540_2 ( .OUT(na2540_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2540_1_i) );
// C_MX2b/D///      x71y65     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2541_1 ( .OUT(na2541_1_i), .IN1(1'b1), .IN2(~na5953_2), .IN3(1'b0), .IN4(1'b0), .IN5(na5249_2), .IN6(na5233_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2541_2 ( .OUT(na2541_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2541_1_i) );
// C_MX2b/D///      x76y57     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2542_1 ( .OUT(na2542_1_i), .IN1(1'b1), .IN2(na5953_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na5234_2), .IN8(na9880_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2542_2 ( .OUT(na2542_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2542_1_i) );
// C_MX2b/D///      x74y64     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2543_1 ( .OUT(na2543_1_i), .IN1(1'b1), .IN2(~na5953_2), .IN3(1'b0), .IN4(1'b0), .IN5(na5251_2), .IN6(na5235_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2543_2 ( .OUT(na2543_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2543_1_i) );
// C_ORAND*/D///      x71y60     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2544_1 ( .OUT(na2544_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9882_2), .IN6(~na5953_2), .IN7(na2521_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2544_2 ( .OUT(na2544_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2544_1_i) );
// C_///ORAND*/D      x63y68     80'h00_F600_80_0000_0C07_FFA7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a2545_4 ( .OUT(na2545_2_i), .IN1(~na5253_2), .IN2(~na5953_2), .IN3(na2523_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2545_5 ( .OUT(na2545_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2545_2_i) );
// C_ORAND*/D///      x71y62     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2546_1 ( .OUT(na2546_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9884_2), .IN6(~na5953_2), .IN7(na2525_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2546_2 ( .OUT(na2546_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2546_1_i) );
// C_///ORAND*/D      x78y68     80'h00_F600_80_0000_0C07_FFC7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a2547_4 ( .OUT(na2547_2_i), .IN1(~na9885_2), .IN2(~na5953_2), .IN3(1'b0), .IN4(na2527_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2547_5 ( .OUT(na2547_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2547_2_i) );
// C_ORAND*/D///      x74y68     80'h00_F600_00_0000_0388_C7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2548_1 ( .OUT(na2548_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9886_2), .IN6(~na5953_2), .IN7(1'b0),
                      .IN8(na2529_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2548_2 ( .OUT(na2548_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2548_1_i) );
// C_ORAND*/D///      x70y72     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2549_1 ( .OUT(na2549_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9887_2), .IN6(~na5953_2), .IN7(na2531_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2549_2 ( .OUT(na2549_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2549_1_i) );
// C_ORAND*/D///      x76y69     80'h00_F600_00_0000_0388_A7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a2550_1 ( .OUT(na2550_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9888_2), .IN6(~na5953_2), .IN7(na2533_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2550_2 ( .OUT(na2550_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2550_1_i) );
// C_///ORAND*/D      x76y69     80'h00_F600_80_0000_0C07_FFA7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a2551_4 ( .OUT(na2551_2_i), .IN1(~na5259_2), .IN2(~na5953_2), .IN3(na2535_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2551_5 ( .OUT(na2551_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2551_2_i) );
// C_MX2b/D///      x76y73     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2552_1 ( .OUT(na2552_1_i), .IN1(1'b1), .IN2(na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1904_1), .IN8(na6014_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2552_2 ( .OUT(na2552_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2552_1_i) );
// C_MX2b/D///      x75y70     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2553_1 ( .OUT(na2553_1_i), .IN1(1'b1), .IN2(na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1922_1), .IN8(na6015_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2553_2 ( .OUT(na2553_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2553_1_i) );
// C_MX2b/D///      x73y80     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2554_1 ( .OUT(na2554_1_i), .IN1(1'b1), .IN2(na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1932_1), .IN8(na6016_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2554_2 ( .OUT(na2554_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2554_1_i) );
// C_MX2b/D///      x75y69     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2555_1 ( .OUT(na2555_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6017_1), .IN8(na1942_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2555_2 ( .OUT(na2555_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2555_1_i) );
// C_MX2b/D///      x72y78     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2556_1 ( .OUT(na2556_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6018_2), .IN6(na1951_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2556_2 ( .OUT(na2556_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2556_1_i) );
// C_MX2b/D///      x75y76     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2557_1 ( .OUT(na2557_1_i), .IN1(1'b1), .IN2(na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1960_1), .IN6(na6019_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2557_2 ( .OUT(na2557_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2557_1_i) );
// C_MX2b/D///      x76y61     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2558_1 ( .OUT(na2558_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6020_2), .IN6(na1969_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2558_2 ( .OUT(na2558_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2558_1_i) );
// C_MX2b/D///      x75y71     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2559_1 ( .OUT(na2559_1_i), .IN1(1'b1), .IN2(na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1978_1), .IN6(na6021_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2559_2 ( .OUT(na2559_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2559_1_i) );
// C_MX2b/D///      x78y71     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2560_1 ( .OUT(na2560_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6022_2), .IN8(na1987_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2560_2 ( .OUT(na2560_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2560_1_i) );
// C_MX2b/D///      x79y72     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2561_1 ( .OUT(na2561_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6023_1), .IN8(na1994_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2561_2 ( .OUT(na2561_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2561_1_i) );
// C_MX2b/D///      x75y77     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2562_1 ( .OUT(na2562_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6024_2), .IN8(na2001_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2562_2 ( .OUT(na2562_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2562_1_i) );
// C_MX2b/D///      x78y76     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2563_1 ( .OUT(na2563_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(na6025_1), .IN6(na2008_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2563_2 ( .OUT(na2563_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2563_1_i) );
// C_MX2b/D///      x71y78     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2564_1 ( .OUT(na2564_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6026_2), .IN8(na2015_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2564_2 ( .OUT(na2564_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2564_1_i) );
// C_MX2b/D///      x71y79     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2565_1 ( .OUT(na2565_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na9212_2), .IN5(1'b0), .IN6(na6027_1), .IN7(1'b0), .IN8(na2022_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2565_2 ( .OUT(na2565_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2565_1_i) );
// C_MX2b/D///      x75y67     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2566_1 ( .OUT(na2566_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6028_2), .IN8(na2029_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2566_2 ( .OUT(na2566_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2566_1_i) );
// C_MX2b/D///      x79y74     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2567_1 ( .OUT(na2567_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6039_1), .IN8(na2106_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2567_2 ( .OUT(na2567_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2567_1_i) );
// C_MX2b/D///      x72y77     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2568_1 ( .OUT(na2568_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6040_2), .IN8(na2113_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2568_2 ( .OUT(na2568_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2568_1_i) );
// C_MX2b/D///      x75y79     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2569_1 ( .OUT(na2569_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6041_1), .IN8(na2120_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2569_2 ( .OUT(na2569_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2569_1_i) );
// C_MX2b/D///      x73y77     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2570_1 ( .OUT(na2570_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6042_2), .IN8(na2127_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2570_2 ( .OUT(na2570_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2570_1_i) );
// C_MX2b/D///      x79y80     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2571_1 ( .OUT(na2571_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6043_1), .IN8(na2134_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2571_2 ( .OUT(na2571_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2571_1_i) );
// C_MX2b/D///      x76y80     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2572_1 ( .OUT(na2572_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6044_2), .IN8(na2141_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2572_2 ( .OUT(na2572_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2572_1_i) );
// C_MX2b/D///      x74y78     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2573_1 ( .OUT(na2573_1_i), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6045_1), .IN8(na2148_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2573_2 ( .OUT(na2573_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2573_1_i) );
// C_MX2b////D      x67y55     80'h00_FE18_00_0040_0A32_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2574_1 ( .OUT(na2574_1), .IN1(1'b1), .IN2(~na343_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2574_2), .IN6(~na2575_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2574_5 ( .OUT(na2574_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2574_1) );
// C_MX2b////      x75y68     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2575_1 ( .OUT(na2575_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6029_1), .IN6(~na2036_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x67y51     80'h00_FE18_00_0040_0A32_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2576_1 ( .OUT(na2576_1), .IN1(1'b1), .IN2(~na343_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2576_2), .IN6(~na2577_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2576_5 ( .OUT(na2576_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2576_1) );
// C_MX2b////      x75y72     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2577_1 ( .OUT(na2577_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6030_2), .IN6(~na2043_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x61y50     80'h00_FE18_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2578_1 ( .OUT(na2578_1), .IN1(1'b1), .IN2(na343_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2579_1), .IN6(na2578_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2578_5 ( .OUT(na2578_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2578_1) );
// C_MX2b////      x75y65     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2579_1 ( .OUT(na2579_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6031_1), .IN6(~na2050_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x70y56     80'h00_FE18_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2580_1 ( .OUT(na2580_1), .IN1(1'b1), .IN2(na343_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2581_1), .IN8(na2580_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2580_5 ( .OUT(na2580_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2580_1) );
// C_MX2b////      x106y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2581_1 ( .OUT(na2581_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6032_2), .IN6(~na2057_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x62y52     80'h00_FE18_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2582_1 ( .OUT(na2582_1), .IN1(1'b1), .IN2(na343_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2583_1), .IN8(na2582_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2582_5 ( .OUT(na2582_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2582_1) );
// C_MX2b////      x82y75     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2583_1 ( .OUT(na2583_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na6033_1), .IN8(~na2064_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x75y85     80'h00_FE18_00_0040_0A32_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2584_1 ( .OUT(na2584_1), .IN1(1'b1), .IN2(~na343_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2584_2), .IN6(~na2585_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2584_5 ( .OUT(na2584_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2584_1) );
// C_MX2b////      x81y74     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2585_1 ( .OUT(na2585_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6034_2), .IN6(~na2071_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x75y96     80'h00_FE18_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2586_1 ( .OUT(na2586_1), .IN1(1'b1), .IN2(na343_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2587_1), .IN6(na2586_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2586_5 ( .OUT(na2586_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2586_1) );
// C_MX2b////      x79y75     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2587_1 ( .OUT(na2587_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na6035_1), .IN8(~na2078_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x76y79     80'h00_FE18_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2588_1 ( .OUT(na2588_1), .IN1(1'b1), .IN2(~na343_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2588_2), .IN8(~na2589_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2588_5 ( .OUT(na2588_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2588_1) );
// C_MX2b////      x54y78     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2589_1 ( .OUT(na2589_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6036_2), .IN6(~na2085_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x76y78     80'h00_FE18_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2590_1 ( .OUT(na2590_1), .IN1(1'b1), .IN2(na343_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2591_1), .IN8(na2590_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2590_5 ( .OUT(na2590_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2590_1) );
// C_MX2b////      x82y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2591_1 ( .OUT(na2591_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na6037_1), .IN6(~na2092_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x76y62     80'h00_FE18_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2592_1 ( .OUT(na2592_1), .IN1(1'b1), .IN2(na343_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2593_1), .IN8(na2592_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2592_5 ( .OUT(na2592_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2592_1) );
// C_MX2b////      x84y77     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2593_1 ( .OUT(na2593_1), .IN1(1'b1), .IN2(~na401_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na6038_2), .IN8(~na2099_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x61y80     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2594_1 ( .OUT(na2594_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na528_1), .IN6(1'b0), .IN7(na6530_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2594_2 ( .OUT(na2594_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2594_1_i) );
// C_MX2b////      x57y83     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2595_1 ( .OUT(na2595_1), .IN1(1'b1), .IN2(na9500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na357_1), .IN8(na9632_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x74y93     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2596_1 ( .OUT(na2596_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na533_1), .IN6(1'b0), .IN7(na6531_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2596_2 ( .OUT(na2596_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2596_1_i) );
// C_MX2b/D///      x70y87     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2597_1 ( .OUT(na2597_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na537_1), .IN6(1'b0), .IN7(na6532_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2597_2 ( .OUT(na2597_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2597_1_i) );
// C_MX2b/D///      x70y91     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2598_1 ( .OUT(na2598_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6533_1), .IN7(1'b0), .IN8(~na3539_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2598_2 ( .OUT(na2598_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2598_1_i) );
// C_MX2b/D///      x65y87     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2599_1 ( .OUT(na2599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6534_1), .IN7(1'b0), .IN8(~na548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2599_2 ( .OUT(na2599_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2599_1_i) );
// C_MX2b/D///      x70y89     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2600_1 ( .OUT(na2600_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6535_1), .IN7(1'b0), .IN8(~na555_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2600_2 ( .OUT(na2600_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2600_1_i) );
// C_MX2b/D///      x68y89     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2601_1 ( .OUT(na2601_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6536_1), .IN7(1'b0), .IN8(~na576_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2601_2 ( .OUT(na2601_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2601_1_i) );
// C_MX2b/D///      x68y82     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2602_1 ( .OUT(na2602_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6537_1), .IN7(1'b0), .IN8(~na584_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2602_2 ( .OUT(na2602_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2602_1_i) );
// C_MX2b/D///      x71y86     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2603_1 ( .OUT(na2603_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na590_1), .IN6(1'b0), .IN7(na6538_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2603_2 ( .OUT(na2603_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2603_1_i) );
// C_MX2b/D///      x70y81     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2604_1 ( .OUT(na2604_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6539_1), .IN7(1'b0), .IN8(~na595_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2604_2 ( .OUT(na2604_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2604_1_i) );
// C_MX2b/D///      x67y87     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2605_1 ( .OUT(na2605_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6540_1), .IN7(1'b0), .IN8(~na600_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2605_2 ( .OUT(na2605_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2605_1_i) );
// C_MX2b/D///      x65y91     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2606_1 ( .OUT(na2606_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6541_1), .IN7(1'b0), .IN8(~na1395_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2606_2 ( .OUT(na2606_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2606_1_i) );
// C_MX2b/D///      x66y96     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2607_1 ( .OUT(na2607_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6542_1), .IN7(1'b0), .IN8(~na604_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2607_2 ( .OUT(na2607_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2607_1_i) );
// C_MX2b/D///      x61y92     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2608_1 ( .OUT(na2608_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6543_1), .IN7(1'b0), .IN8(~na610_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2608_2 ( .OUT(na2608_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2608_1_i) );
// C_MX2b/D///      x70y94     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2609_1 ( .OUT(na2609_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na620_1), .IN6(1'b0), .IN7(na6544_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2609_2 ( .OUT(na2609_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2609_1_i) );
// C_MX2b/D///      x66y83     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2610_1 ( .OUT(na2610_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6545_1), .IN7(1'b0), .IN8(~na615_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2610_2 ( .OUT(na2610_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2610_1_i) );
// C_MX2b/D///      x74y92     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2611_1 ( .OUT(na2611_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6546_1), .IN7(1'b0), .IN8(~na625_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2611_2 ( .OUT(na2611_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2611_1_i) );
// C_MX2b/D///      x66y85     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2612_1 ( .OUT(na2612_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na1601_1), .IN6(1'b0), .IN7(na6547_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2612_2 ( .OUT(na2612_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2612_1_i) );
// C_MX2b/D///      x66y91     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2613_1 ( .OUT(na2613_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6548_1), .IN7(1'b0), .IN8(~na630_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2613_2 ( .OUT(na2613_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2613_1_i) );
// C_MX2b/D///      x66y90     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2614_1 ( .OUT(na2614_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6549_1), .IN7(1'b0), .IN8(~na635_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2614_2 ( .OUT(na2614_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2614_1_i) );
// C_MX2b/D///      x68y96     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2615_1 ( .OUT(na2615_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na1584_1), .IN6(1'b0), .IN7(na6550_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2615_2 ( .OUT(na2615_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2615_1_i) );
// C_MX2b/D///      x68y91     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2616_1 ( .OUT(na2616_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6551_1), .IN7(1'b0), .IN8(~na659_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2616_2 ( .OUT(na2616_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2616_1_i) );
// C_MX2b/D///      x73y96     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2617_1 ( .OUT(na2617_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6552_1), .IN7(1'b0), .IN8(~na665_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2617_2 ( .OUT(na2617_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2617_1_i) );
// C_MX2b/D///      x61y93     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2618_1 ( .OUT(na2618_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6553_1), .IN7(1'b0), .IN8(~na670_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2618_2 ( .OUT(na2618_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2618_1_i) );
// C_MX2b/D///      x73y95     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2619_1 ( .OUT(na2619_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6554_1), .IN7(1'b0), .IN8(~na675_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2619_2 ( .OUT(na2619_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2619_1_i) );
// C_MX2b/D///      x72y95     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2620_1 ( .OUT(na2620_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6555_1), .IN7(1'b0), .IN8(~na680_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2620_2 ( .OUT(na2620_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2620_1_i) );
// C_MX2b/D///      x69y96     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2621_1 ( .OUT(na2621_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na685_1), .IN6(1'b0), .IN7(na6556_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2621_2 ( .OUT(na2621_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2621_1_i) );
// C_MX2b/D///      x65y95     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2622_1 ( .OUT(na2622_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6557_1), .IN7(1'b0), .IN8(~na690_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2622_2 ( .OUT(na2622_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2622_1_i) );
// C_MX2b/D///      x68y101     80'h00_F600_00_0040_0A51_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2623_1 ( .OUT(na2623_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na359_1), .IN4(1'b1), .IN5(~na695_1), .IN6(1'b0), .IN7(na6558_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2623_2 ( .OUT(na2623_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2623_1_i) );
// C_MX2b/D///      x74y95     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2624_1 ( .OUT(na2624_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6559_1), .IN7(1'b0), .IN8(~na700_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2624_2 ( .OUT(na2624_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2624_1_i) );
// C_MX2b/D///      x67y93     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2625_1 ( .OUT(na2625_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6560_1), .IN7(1'b0), .IN8(~na705_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2625_2 ( .OUT(na2625_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2625_1_i) );
// C_MX2b/D///      x65y94     80'h00_F600_00_0040_0AA8_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2626_1 ( .OUT(na2626_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na359_1), .IN4(1'b1), .IN5(1'b0), .IN6(na6561_1), .IN7(1'b0), .IN8(~na720_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2626_2 ( .OUT(na2626_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2626_1_i) );
// C_XOR////      x54y59     80'h00_0018_02_0800_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2627_1 ( .OUT(na2627_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na50_1), .IN6(na3598_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_2080)) 
           _a2627_6 ( .COUTY1(na2627_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na2627_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX4b/D///      x117y122     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2659_1 ( .OUT(na2659_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1081_1), .IN6(~na2660_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2659_2 ( .OUT(na2659_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2659_1_i) );
// C_MX2b////      x111y96     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2660_1 ( .OUT(na2660_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1275_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na3992_2), .IN7(1'b0), .IN8(~na1161_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x122y96     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2661_1 ( .OUT(na2661_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9648_2), .IN6(na454_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2661_2 ( .OUT(na2661_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2661_1_i) );
// C_MX4b/D///      x116y119     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2662_1 ( .OUT(na2662_1_i), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1075_1), .IN6(~na2663_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2662_2 ( .OUT(na2662_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2662_1_i) );
// C_MX2b////      x113y104     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2663_1 ( .OUT(na2663_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1275_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na4019_2), .IN7(1'b0), .IN8(~na1156_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x113y120     80'h00_FE00_00_0040_0A31_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2664_1 ( .OUT(na2664_1_i), .IN1(~na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na2665_1), .IN6(na1074_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2664_2 ( .OUT(na2664_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2664_1_i) );
// C_MX2b////      x111y123     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2665_1 ( .OUT(na2665_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1275_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na4019_1), .IN7(1'b0), .IN8(~na1155_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x113y114     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2666_1 ( .OUT(na2666_1_i), .IN1(na1215_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9649_2),
                      .IN8(na1289_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2666_2 ( .OUT(na2666_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2666_1_i) );
// C_MX4b/D///      x109y107     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2667_1 ( .OUT(na2667_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2667_1), .IN6(na1211_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2667_2 ( .OUT(na2667_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2667_1_i) );
// C_MX4b/D///      x101y110     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2668_1 ( .OUT(na2668_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1139_1), .IN6(na2668_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2668_2 ( .OUT(na2668_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2668_1_i) );
// C_MX4b/D///      x113y109     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2669_1 ( .OUT(na2669_1_i), .IN1(1'b1), .IN2(na1073_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2669_1), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2669_2 ( .OUT(na2669_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2669_1_i) );
// C_MX4b/D///      x109y103     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2670_1 ( .OUT(na2670_1_i), .IN1(1'b1), .IN2(~na1073_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na9651_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2670_2 ( .OUT(na2670_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2670_1_i) );
// C_MX4b/D///      x113y94     80'h00_FE00_00_0040_0A31_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2671_1 ( .OUT(na2671_1_i), .IN1(1'b1), .IN2(~na996_2), .IN3(1'b1), .IN4(na6626_1), .IN5(~na2672_1), .IN6(na2671_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2671_2 ( .OUT(na2671_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2671_1_i) );
// C_MX2b////      x121y97     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2672_1 ( .OUT(na2672_1), .IN1(1'b0), .IN2(1'b0), .IN3(na997_1), .IN4(1'b1), .IN5(~na3972_1), .IN6(1'b0), .IN7(~na3865_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x116y95     80'h00_FE00_00_0040_0AC8_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2673_1 ( .OUT(na2673_1_i), .IN1(1'b1), .IN2(na996_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2673_1),
                      .IN8(~na9652_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2673_2 ( .OUT(na2673_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2673_1_i) );
// C_AND/D///      x110y91     80'h00_FE00_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2675_1 ( .OUT(na2675_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2676_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2675_2 ( .OUT(na2675_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2675_1_i) );
// C_ANDXOR////      x119y100     80'h00_0018_00_0000_0C66_A700
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a2676_1 ( .OUT(na2676_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na951_1), .IN6(na8058_2), .IN7(~na2675_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x92y93     80'h00_FE00_80_0000_0C88_3335
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2677_1 ( .OUT(na2677_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2678_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2677_2 ( .OUT(na2677_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2677_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2677_4 ( .OUT(na2677_2_i), .IN1(~na1321_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2677_5 ( .OUT(na2677_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2677_2_i) );
// C_MX2a////      x89y88     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2678_1 ( .OUT(na2678_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2677_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1322_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x86y86     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2679_4 ( .OUT(na2679_2_i), .IN1(na2680_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2679_5 ( .OUT(na2679_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2679_2_i) );
// C_AND////      x87y93     80'h00_0018_00_0000_0888_322F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2680_1 ( .OUT(na2680_1), .IN1(1'b1), .IN2(1'b1), .IN3(na436_1), .IN4(~na452_1), .IN5(na428_1), .IN6(~na435_1), .IN7(1'b1),
                      .IN8(~na452_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x100y93     80'h00_FE00_80_0000_0C88_1F33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2681_1 ( .OUT(na2681_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2682_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2681_2 ( .OUT(na2681_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2681_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2681_4 ( .OUT(na2681_2_i), .IN1(1'b1), .IN2(~na1236_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2681_5 ( .OUT(na2681_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2681_2_i) );
// C_MX2a////      x94y87     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2682_1 ( .OUT(na2682_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2681_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na1237_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x85y81     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2684_1 ( .OUT(na2684_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1355_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1357_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x84y85     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2686_1 ( .OUT(na2686_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1359_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na1361_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x78y77     80'h00_FE00_80_0000_0C88_1F33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2687_1 ( .OUT(na2687_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2688_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2687_2 ( .OUT(na2687_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2687_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2687_4 ( .OUT(na2687_2_i), .IN1(1'b1), .IN2(~na2691_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2687_5 ( .OUT(na2687_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2687_2_i) );
// C_MX2a////      x88y87     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2688_1 ( .OUT(na2688_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2687_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na2689_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y84     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2689_4 ( .OUT(na2689_2), .IN1(na566_1), .IN2(~na435_1), .IN3(na433_2), .IN4(na9230_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x85y80     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2691_1 ( .OUT(na2691_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2687_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na2689_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x50y111     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2692_1 ( .OUT(na2692_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3833_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2692_2 ( .OUT(na2692_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2692_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2692_4 ( .OUT(na2692_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(na3833_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2692_5 ( .OUT(na2692_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2692_2_i) );
// C_MX4b/D///      x109y93     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2693_1 ( .OUT(na2693_1_i), .IN1(~na954_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na9659_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2693_2 ( .OUT(na2693_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2693_1_i) );
// C_MX4b/D///      x98y70     80'h00_FE00_00_0040_0AC3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2695_1 ( .OUT(na2695_1_i), .IN1(~na2696_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na260_1),
                      .IN8(na2695_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2695_2 ( .OUT(na2695_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2695_1_i) );
// C_///AND/      x99y69     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2696_4 ( .OUT(na2696_2), .IN1(na9229_2), .IN2(1'b1), .IN3(na1471_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x107y73     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2697_1 ( .OUT(na2697_1_i), .IN1(na2696_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2697_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2697_2 ( .OUT(na2697_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2697_1_i) );
// C_MX4b/D///      x98y63     80'h00_FE00_00_0040_0AC3_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2698_1 ( .OUT(na2698_1_i), .IN1(na2696_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na2698_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2698_2 ( .OUT(na2698_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2698_1_i) );
// C_MX4b/D///      x94y59     80'h00_FE00_00_0040_0AC3_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2699_1 ( .OUT(na2699_1_i), .IN1(na426_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na2699_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2699_2 ( .OUT(na2699_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2699_1_i) );
// C_MX4b/D///      x117y98     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2701_1 ( .OUT(na2701_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9661_2), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2701_2 ( .OUT(na2701_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2701_1_i) );
// C_MX4b/D///      x113y99     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2702_1 ( .OUT(na2702_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2702_1), .IN6(na1078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2702_2 ( .OUT(na2702_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2702_1_i) );
// C_MX4b/D///      x117y109     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2703_1 ( .OUT(na2703_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2703_1), .IN6(na1073_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2703_2 ( .OUT(na2703_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2703_1_i) );
// C_MX4b/D///      x114y97     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2704_1 ( .OUT(na2704_1_i), .IN1(1'b1), .IN2(na454_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na9664_2), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2704_2 ( .OUT(na2704_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2704_1_i) );
// C_MX4b/D///      x116y92     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2705_1 ( .OUT(na2705_1_i), .IN1(1'b1), .IN2(~na454_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na2705_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2705_2 ( .OUT(na2705_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2705_1_i) );
// C_///ORAND/D      x112y92     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2706_4 ( .OUT(na2706_2_i), .IN1(na8061_1), .IN2(na2707_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2706_5 ( .OUT(na2706_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2706_2_i) );
// C_AND////      x109y74     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2707_1 ( .OUT(na2707_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2927_1), .IN7(na298_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x128y74     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2708_1 ( .OUT(na2708_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2709_2), .IN6(na8063_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2708_2 ( .OUT(na2708_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2708_1_i) );
// C_///AND/      x113y75     80'h00_0060_00_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2709_4 ( .OUT(na2709_2), .IN1(na2928_1), .IN2(1'b1), .IN3(na298_1), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x126y74     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2710_1 ( .OUT(na2710_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2711_2), .IN6(na8065_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2710_2 ( .OUT(na2710_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2710_1_i) );
// C_///AND/      x115y87     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2711_4 ( .OUT(na2711_2), .IN1(1'b1), .IN2(na9194_2), .IN3(na2929_1), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x126y76     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2712_1 ( .OUT(na2712_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2713_1), .IN6(na8067_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2712_2 ( .OUT(na2712_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2712_1_i) );
// C_AND////      x127y67     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2713_1 ( .OUT(na2713_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2930_1), .IN6(1'b1), .IN7(na298_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x124y74     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2714_1 ( .OUT(na2714_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8069_1), .IN6(na2715_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2714_2 ( .OUT(na2714_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2714_1_i) );
// C_///AND/      x125y62     80'h00_0060_00_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2715_4 ( .OUT(na2715_2), .IN1(na1828_1), .IN2(1'b1), .IN3(na298_1), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x104y92     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2716_1 ( .OUT(na2716_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1095_2),
                      .IN8(na2716_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2716_2 ( .OUT(na2716_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2716_1_i) );
// C_MX4b/D///      x119y89     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2717_1 ( .OUT(na2717_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2717_1), .IN6(na961_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2717_2 ( .OUT(na2717_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2717_1_i) );
// C_AND/D//AND/D      x127y56     80'h00_FE00_80_0000_0C88_1F53
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2718_1 ( .OUT(na2718_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2248_1), .IN8(~na2719_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2718_2 ( .OUT(na2718_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2718_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2718_4 ( .OUT(na2718_2_i), .IN1(1'b1), .IN2(~na2249_1), .IN3(~na2248_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2718_5 ( .OUT(na2718_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2718_2_i) );
// C_MX2b////      x128y54     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2719_1 ( .OUT(na2719_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na500_2), .IN5(1'b0), .IN6(~na2718_1), .IN7(1'b0), .IN8(~na8070_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x103y99     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2720_1 ( .OUT(na2720_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2720_1), .IN6(na893_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2720_2 ( .OUT(na2720_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2720_1_i) );
// C_MX4b/D///      x101y107     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2721_1 ( .OUT(na2721_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9666_2),
                      .IN8(na3761_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2721_2 ( .OUT(na2721_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2721_1_i) );
// C_MX2b////      x101y116     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2722_1 ( .OUT(na2722_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na6057_1), .IN4(1'b1), .IN5(1'b0), .IN6(na4118_1), .IN7(1'b0), .IN8(na2725_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x112y86     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2723_4 ( .OUT(na2723_2_i), .IN1(na8072_1), .IN2(na2724_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2723_5 ( .OUT(na2723_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2723_2_i) );
// C_AND////      x127y70     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2724_1 ( .OUT(na2724_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na9194_2), .IN7(na1418_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////D      x108y110     80'h00_D518_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2725_1 ( .OUT(na2725_1), .IN1(1'b1), .IN2(na316_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1870_1), .IN6(~na2722_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2725_5 ( .OUT(na2725_2), .CLK(~na4116_1), .EN(~na3239_1), .SR(~na1_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2725_1) );
// C_MX2b/D///      x121y96     80'h00_F900_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2726_1 ( .OUT(na2726_1_i), .IN1(1'b1), .IN2(na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(na935_1), .IN6(na3167_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2726_2 ( .OUT(na2726_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2726_1_i) );
// C_MX2b/D///      x112y103     80'h00_F900_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2727_1 ( .OUT(na2727_1_i), .IN1(1'b1), .IN2(na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(na936_1), .IN6(na2726_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2727_2 ( .OUT(na2727_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2727_1_i) );
// C_MX2b/D///      x119y104     80'h00_F900_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2728_1 ( .OUT(na2728_1_i), .IN1(1'b1), .IN2(~na6065_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2727_1), .IN8(na937_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2728_2 ( .OUT(na2728_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2728_1_i) );
// C_MX2b/D///      x124y113     80'h00_F900_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2729_1 ( .OUT(na2729_1_i), .IN1(1'b1), .IN2(na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(na938_1), .IN6(na2728_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2729_2 ( .OUT(na2729_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2729_1_i) );
// C_MX2b/D///      x124y117     80'h00_F900_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2730_1 ( .OUT(na2730_1_i), .IN1(1'b1), .IN2(~na6065_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2729_1), .IN8(na939_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2730_2 ( .OUT(na2730_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2730_1_i) );
// C_MX2b/D///      x123y118     80'h00_F900_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2731_1 ( .OUT(na2731_1_i), .IN1(1'b1), .IN2(~na6065_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2730_1), .IN8(na940_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2731_2 ( .OUT(na2731_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2731_1_i) );
// C_MX2b/D///      x96y90     80'h00_F900_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2732_1 ( .OUT(na2732_1_i), .IN1(1'b1), .IN2(na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(na941_1), .IN6(na2731_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2732_2 ( .OUT(na2732_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2732_1_i) );
// C_MX2b/D///      x113y101     80'h00_F900_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2733_1 ( .OUT(na2733_1_i), .IN1(1'b1), .IN2(na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2693_1), .IN6(~na9667_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2733_2 ( .OUT(na2733_1), .CLK(~na4116_1), .EN(na3238_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2733_1_i) );
// C_OR////DST      x112y100     80'h20_7D18_00_0000_0EEE_AC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2734_1 ( .OUT(na2734_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na316_1), .IN7(na8073_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0000)) 
           _a2734_5 ( .OUT(na2734_2), .CLK(~na4116_1), .EN(1'b1), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2734_1) );
// C_///ORAND/D      x126y57     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2735_4 ( .OUT(na2735_2_i), .IN1(na8075_2), .IN2(na2736_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2735_5 ( .OUT(na2735_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2735_2_i) );
// C_///AND/      x127y58     80'h00_0060_00_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2736_4 ( .OUT(na2736_2), .IN1(na3191_1), .IN2(1'b1), .IN3(na298_1), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x126y55     80'h00_FE00_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2737_1 ( .OUT(na2737_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2248_1), .IN8(~na2738_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2737_2 ( .OUT(na2737_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2737_1_i) );
// C_MX2b////      x130y52     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2738_1 ( .OUT(na2738_1), .IN1(1'b1), .IN2(na9244_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2737_1), .IN8(~na8076_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x102y108     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2739_1 ( .OUT(na2739_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3759_1),
                      .IN8(na2739_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2739_2 ( .OUT(na2739_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2739_1_i) );
// C_MX4b/D///      x112y95     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2740_1 ( .OUT(na2740_1_i), .IN1(na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9668_2), .IN6(na1073_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2740_2 ( .OUT(na2740_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2740_1_i) );
// C_MX4b/D///      x113y93     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2741_1 ( .OUT(na2741_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2741_1), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2741_2 ( .OUT(na2741_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2741_1_i) );
// C_MX4b/D///      x107y81     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2743_1 ( .OUT(na2743_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2743_1), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2743_2 ( .OUT(na2743_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2743_1_i) );
// C_MX4b/D///      x105y105     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2744_1 ( .OUT(na2744_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2744_1), .IN6(na1078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2744_2 ( .OUT(na2744_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2744_1_i) );
// C_MX4b/D///      x119y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2745_1 ( .OUT(na2745_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2745_1), .IN6(na1091_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2745_2 ( .OUT(na2745_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2745_1_i) );
// C_///AND/D      x127y57     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2746_4 ( .OUT(na2746_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na2248_1), .IN4(~na2747_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2746_5 ( .OUT(na2746_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2746_2_i) );
// C_MX2b////      x126y52     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2747_1 ( .OUT(na2747_1), .IN1(1'b1), .IN2(na9244_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2746_2), .IN6(~na8077_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x96y107     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2748_1 ( .OUT(na2748_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2748_1),
                      .IN8(na3761_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2748_2 ( .OUT(na2748_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2748_1_i) );
// C_MX2b////      x75y36     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2749_1 ( .OUT(na2749_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na6058_2), .IN4(1'b1), .IN5(na4119_2), .IN6(1'b0), .IN7(na2751_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x112y84     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2750_1 ( .OUT(na2750_1_i), .IN1(1'b1), .IN2(~na1160_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na2750_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2750_2 ( .OUT(na2750_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2750_1_i) );
// C_MX2b////D      x88y43     80'h00_D518_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2751_1 ( .OUT(na2751_1), .IN1(1'b1), .IN2(na9506_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2833_1), .IN6(~na2749_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2751_5 ( .OUT(na2751_2), .CLK(~na4116_1), .EN(~na3275_1), .SR(~na2_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2751_1) );
// C_MX2b/D///      x106y67     80'h00_F900_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2752_1 ( .OUT(na2752_1_i), .IN1(na6118_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2828_1), .IN6(na1419_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2752_2 ( .OUT(na2752_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2752_1_i) );
// C_MX2b/D///      x108y67     80'h00_F900_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2753_1 ( .OUT(na2753_1_i), .IN1(~na6118_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2752_1), .IN8(na2827_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2753_2 ( .OUT(na2753_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2753_1_i) );
// C_MX2b/D///      x105y68     80'h00_F900_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2754_1 ( .OUT(na2754_1_i), .IN1(~na6118_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2753_1), .IN8(na2826_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2754_2 ( .OUT(na2754_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2754_1_i) );
// C_MX2b/D///      x112y71     80'h00_F900_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2755_1 ( .OUT(na2755_1_i), .IN1(na6118_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2825_1), .IN6(na2754_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2755_2 ( .OUT(na2755_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2755_1_i) );
// C_MX2b/D///      x104y71     80'h00_F900_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2756_1 ( .OUT(na2756_1_i), .IN1(~na6118_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2755_1), .IN8(na2824_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2756_2 ( .OUT(na2756_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2756_1_i) );
// C_MX2b/D///      x103y70     80'h00_F900_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2757_1 ( .OUT(na2757_1_i), .IN1(~na6118_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2756_1), .IN8(na2823_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2757_2 ( .OUT(na2757_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2757_1_i) );
// C_MX2b/D///      x93y61     80'h00_F900_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2758_1 ( .OUT(na2758_1_i), .IN1(na6118_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2821_1), .IN6(na2757_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2758_2 ( .OUT(na2758_1), .CLK(~na4116_1), .EN(na3255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2758_1_i) );
// C_MX2b/D///      x109y66     80'h00_F900_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2759_1 ( .OUT(na2759_1_i), .IN1(na6118_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2832_1), .IN6(~na2759_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2759_2 ( .OUT(na2759_1), .CLK(~na4116_1), .EN(na3254_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2759_1_i) );
// C_OR////DST      x107y66     80'h20_7D18_00_0000_0EEE_E000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a2760_1 ( .OUT(na2760_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8078_1), .IN8(na1425_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0000)) 
           _a2760_5 ( .OUT(na2760_2), .CLK(~na4116_1), .EN(1'b1), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2760_1) );
// C_MX4b/D///      x106y104     80'h00_FE00_00_0040_0AC3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2761_1 ( .OUT(na2761_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na833_1),
                      .IN8(na2761_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2761_2 ( .OUT(na2761_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2761_1_i) );
// C_MX4b/D///      x120y95     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2762_1 ( .OUT(na2762_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9672_2), .IN6(na1078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2762_2 ( .OUT(na2762_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2762_1_i) );
// C_AND////      x99y64     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2763_1 ( .OUT(na2763_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9947_2), .IN6(1'b1), .IN7(1'b1), .IN8(na6673_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x113y83     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2764_1 ( .OUT(na2764_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2764_1), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2764_2 ( .OUT(na2764_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2764_1_i) );
// C_MX2a////      x105y70     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2766_1 ( .OUT(na2766_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2811_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na2767_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y84     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2767_1 ( .OUT(na2767_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9954_2), .IN6(~na435_1), .IN7(na436_1), .IN8(~na452_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x129y74     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2768_4 ( .OUT(na2768_2_i), .IN1(na8080_1), .IN2(na2772_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2768_5 ( .OUT(na2768_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2768_2_i) );
// C_///AND/      x129y70     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2769_4 ( .OUT(na2769_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na2770_1), .IN4(na8081_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y75     80'h00_0018_00_0000_0888_7F7C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2770_1 ( .OUT(na2770_1), .IN1(1'b0), .IN2(na99_2), .IN3(~na2788_1), .IN4(~na1036_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na2787_1),
                      .IN8(~na1036_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y73     80'h00_0018_00_0000_0C88_7CFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2771_1 ( .OUT(na2771_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na99_2), .IN7(~na2787_1), .IN8(~na1036_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x127y74     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2772_4 ( .OUT(na2772_2), .IN1(1'b1), .IN2(na99_2), .IN3(na2787_1), .IN4(na1036_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x79y78     80'h00_FE00_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2773_1 ( .OUT(na2773_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na8085_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2773_2 ( .OUT(na2773_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2773_1_i) );
// C_ORAND/D///      x122y74     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2774_1 ( .OUT(na2774_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2775_1), .IN6(na8087_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2774_2 ( .OUT(na2774_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2774_1_i) );
// C_AND////      x129y67     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2775_1 ( .OUT(na2775_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na443_1), .IN6(1'b1), .IN7(na298_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x120y68     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2776_1 ( .OUT(na2776_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2777_2), .IN6(na8089_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2776_2 ( .OUT(na2776_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2776_1_i) );
// C_///AND/      x127y59     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2777_4 ( .OUT(na2777_2), .IN1(1'b1), .IN2(na641_1), .IN3(na298_1), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x124y76     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2778_1 ( .OUT(na2778_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2779_1), .IN6(na8091_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2778_2 ( .OUT(na2778_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2778_1_i) );
// C_AND////      x129y69     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2779_1 ( .OUT(na2779_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1653_1), .IN6(1'b1), .IN7(na298_1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x111y94     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2780_1 ( .OUT(na2780_1_i), .IN1(~na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na2780_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2780_2 ( .OUT(na2780_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2780_1_i) );
// C_MX4b/D///      x105y76     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2781_1 ( .OUT(na2781_1_i), .IN1(na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9676_2), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2781_2 ( .OUT(na2781_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2781_1_i) );
// C_MX4b/D///      x111y80     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2782_1 ( .OUT(na2782_1_i), .IN1(~na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na9677_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2782_2 ( .OUT(na2782_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2782_1_i) );
// C_MX4b/D///      x109y72     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2783_1 ( .OUT(na2783_1_i), .IN1(~na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na9678_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2783_2 ( .OUT(na2783_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2783_1_i) );
// C_MX4b/D///      x111y78     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2784_1 ( .OUT(na2784_1_i), .IN1(na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9679_2), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2784_2 ( .OUT(na2784_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2784_1_i) );
// C_MX4b/D///      x104y74     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2785_1 ( .OUT(na2785_1_i), .IN1(~na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na2785_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2785_2 ( .OUT(na2785_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2785_1_i) );
// C_MX4b/D///      x119y76     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2786_1 ( .OUT(na2786_1_i), .IN1(~na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na9680_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2786_2 ( .OUT(na2786_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2786_1_i) );
// C_MX4b/D///      x116y79     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2787_1 ( .OUT(na2787_1_i), .IN1(na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2787_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2787_2 ( .OUT(na2787_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2787_1_i) );
// C_MX4b/D///      x118y77     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2788_1 ( .OUT(na2788_1_i), .IN1(na1037_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9681_2), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2788_2 ( .OUT(na2788_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2788_1_i) );
// C_AND/D//AND*/D      x98y98     80'h00_FE00_80_0000_0C87_3C8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2789_1 ( .OUT(na2789_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1160_2), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2789_2 ( .OUT(na2789_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2789_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a2789_4 ( .OUT(na2789_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2804_1), .IN4(na2789_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2789_5 ( .OUT(na2789_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2789_2_i) );
// C_MX4b/D///      x113y95     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2790_1 ( .OUT(na2790_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2790_1), .IN6(na482_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2790_2 ( .OUT(na2790_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2790_1_i) );
// C_MX4b/D///      x114y94     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2791_1 ( .OUT(na2791_1_i), .IN1(1'b1), .IN2(~na1160_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na833_1),
                      .IN8(na2791_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2791_2 ( .OUT(na2791_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2791_1_i) );
// C_MX4b/D///      x117y105     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2792_1 ( .OUT(na2792_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2792_1), .IN6(na893_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2792_2 ( .OUT(na2792_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2792_1_i) );
// C_MX4b/D///      x123y101     80'h00_FE00_00_0040_0A3C_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2793_1 ( .OUT(na2793_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2793_1), .IN6(na454_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2793_2 ( .OUT(na2793_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2793_1_i) );
// C_MX4b/D///      x121y103     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2794_1 ( .OUT(na2794_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2794_1), .IN6(na1078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2794_2 ( .OUT(na2794_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2794_1_i) );
// C_MX4b/D///      x119y112     80'h00_FE00_00_0040_0A3C_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2795_1 ( .OUT(na2795_1_i), .IN1(1'b1), .IN2(~na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na2795_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2795_2 ( .OUT(na2795_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2795_1_i) );
// C_MX4b/D///      x117y111     80'h00_FE00_00_0040_0A3C_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2796_1 ( .OUT(na2796_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2796_1), .IN6(na1073_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2796_2 ( .OUT(na2796_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2796_1_i) );
// C_MX4b/D///      x95y103     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2797_1 ( .OUT(na2797_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2797_1), .IN6(na1103_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2797_2 ( .OUT(na2797_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2797_1_i) );
// C_MX4b/D///      x112y80     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2798_1 ( .OUT(na2798_1_i), .IN1(1'b1), .IN2(~na1160_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na2798_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2798_2 ( .OUT(na2798_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2798_1_i) );
// C_MX2b////      x125y51     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2800_1 ( .OUT(na2800_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na500_2), .IN5(~na985_2), .IN6(1'b0), .IN7(~na8092_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x108y78     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2801_1 ( .OUT(na2801_1_i), .IN1(1'b1), .IN2(~na1160_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na2801_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2801_2 ( .OUT(na2801_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2801_1_i) );
// C_MX4b/D///      x119y83     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2802_1 ( .OUT(na2802_1_i), .IN1(1'b1), .IN2(~na1160_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na9686_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2802_2 ( .OUT(na2802_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2802_1_i) );
// C_MX4b/D///      x111y83     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2803_1 ( .OUT(na2803_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2803_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2803_2 ( .OUT(na2803_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2803_1_i) );
// C_MX4b/D///      x102y103     80'h00_FE00_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2804_1 ( .OUT(na2804_1_i), .IN1(1'b1), .IN2(na1160_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2804_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2804_2 ( .OUT(na2804_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2804_1_i) );
// C_AND/D//AND/D      x120y81     80'h00_FE00_80_0000_0C88_1F33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2805_1 ( .OUT(na2805_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2806_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2805_2 ( .OUT(na2805_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2805_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2805_4 ( .OUT(na2805_2_i), .IN1(1'b1), .IN2(~na2817_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2805_5 ( .OUT(na2805_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2805_2_i) );
// C_MX2a////      x104y83     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2806_1 ( .OUT(na2806_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2805_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na2807_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y84     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2807_4 ( .OUT(na2807_2), .IN1(~na9226_2), .IN2(na435_2), .IN3(na436_1), .IN4(~na452_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x106y71     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2808_4 ( .OUT(na2808_2_i), .IN1(na2809_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2808_5 ( .OUT(na2808_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2808_2_i) );
// C_AND////      x101y73     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2809_1 ( .OUT(na2809_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na955_1), .IN7(na2810_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y79     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2810_1 ( .OUT(na2810_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9229_2), .IN6(~na435_1), .IN7(na433_2), .IN8(~na452_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x118y83     80'h00_FE00_80_0000_0C88_1F33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2811_1 ( .OUT(na2811_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2812_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2811_2 ( .OUT(na2811_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2811_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2811_4 ( .OUT(na2811_2_i), .IN1(1'b1), .IN2(~na2766_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2811_5 ( .OUT(na2811_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2811_2_i) );
// C_MX2a////      x104y91     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2812_1 ( .OUT(na2812_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2811_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na2767_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x123y87     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2814_1 ( .OUT(na2814_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2818_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na2815_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y94     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2815_1 ( .OUT(na2815_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9229_2), .IN6(~na435_1), .IN7(na433_1), .IN8(~na452_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x109y76     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2817_1 ( .OUT(na2817_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2805_2), .IN4(~na159_1), .IN5(na428_1), .IN6(na2807_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x112y83     80'h00_FE00_80_0000_0C88_1F35
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2818_1 ( .OUT(na2818_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2819_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2818_2 ( .OUT(na2818_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2818_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2818_4 ( .OUT(na2818_2_i), .IN1(~na2814_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2818_5 ( .OUT(na2818_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2818_2_i) );
// C_MX2a////      x102y87     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2819_1 ( .OUT(na2819_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2818_1), .IN4(~na159_1), .IN5(na853_2), .IN6(na2815_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x122y76     80'h00_FE00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2820_1 ( .OUT(na2820_1_i), .IN1(1'b1), .IN2(~na2769_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2771_1),
                      .IN8(na2820_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2820_2 ( .OUT(na2820_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2820_1_i) );
// C_MX4b/D///      x107y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2821_1 ( .OUT(na2821_1_i), .IN1(na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2821_1), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2821_2 ( .OUT(na2821_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2821_1_i) );
// C_AND////      x111y65     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2822_1 ( .OUT(na2822_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(1'b1), .IN7(na2810_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x114y64     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2823_1 ( .OUT(na2823_1_i), .IN1(~na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na2823_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2823_2 ( .OUT(na2823_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2823_1_i) );
// C_MX4b/D///      x114y68     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2824_1 ( .OUT(na2824_1_i), .IN1(~na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na2824_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2824_2 ( .OUT(na2824_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2824_1_i) );
// C_MX4b/D///      x113y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2825_1 ( .OUT(na2825_1_i), .IN1(na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2825_1), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2825_2 ( .OUT(na2825_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2825_1_i) );
// C_MX4b/D///      x120y70     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2826_1 ( .OUT(na2826_1_i), .IN1(~na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na2826_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2826_2 ( .OUT(na2826_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2826_1_i) );
// C_MX4b/D///      x118y66     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2827_1 ( .OUT(na2827_1_i), .IN1(~na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na2827_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2827_2 ( .OUT(na2827_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2827_1_i) );
// C_MX4b/D///      x115y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2828_1 ( .OUT(na2828_1_i), .IN1(na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2828_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2828_2 ( .OUT(na2828_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2828_1_i) );
// C_MX4b/D///      x112y70     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2829_1 ( .OUT(na2829_1_i), .IN1(na2822_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9694_2),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2829_2 ( .OUT(na2829_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2829_1_i) );
// C_MX4b/D///      x86y63     80'h00_FE00_00_0040_0AC3_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2830_1 ( .OUT(na2830_1_i), .IN1(1'b1), .IN2(na2831_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na2830_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2830_2 ( .OUT(na2830_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2830_1_i) );
// C_///AND/      x99y74     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2831_4 ( .OUT(na2831_2), .IN1(na488_1), .IN2(1'b1), .IN3(na2810_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x109y67     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2832_1 ( .OUT(na2832_1_i), .IN1(~na2809_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na9695_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2832_2 ( .OUT(na2832_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2832_1_i) );
// C_MX4b/D///      x101y63     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2833_1 ( .OUT(na2833_1_i), .IN1(na2809_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2833_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2833_2 ( .OUT(na2833_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2833_1_i) );
// C_MX4b/D///      x109y70     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2834_1 ( .OUT(na2834_1_i), .IN1(na2809_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9696_2),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2834_2 ( .OUT(na2834_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2834_1_i) );
// C_AND/D//AND/D      x101y79     80'h00_FE00_80_0000_0C88_2824
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2835_1 ( .OUT(na2835_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na428_2), .IN6(na435_1), .IN7(na433_2), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2835_2 ( .OUT(na2835_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2835_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2835_4 ( .OUT(na2835_2_i), .IN1(~na7072_1), .IN2(na435_1), .IN3(na433_1), .IN4(~na452_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2835_5 ( .OUT(na2835_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2835_2_i) );
// C_///AND/D      x108y90     80'h00_FE00_80_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2836_4 ( .OUT(na2836_2_i), .IN1(1'b1), .IN2(~na8093_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2836_5 ( .OUT(na2836_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2836_2_i) );
// C_AND/D///      x112y81     80'h00_FE00_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2838_1 ( .OUT(na2838_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3542_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2838_2 ( .OUT(na2838_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2838_1_i) );
// C_AND////      x65y93     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2839_1 ( .OUT(na2839_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2843_1), .IN8(na2840_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x72y68     80'h00_0018_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2840_1 ( .OUT(na2840_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na155_1), .IN6(na8095_1), .IN7(1'b0), .IN8(na2841_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y70     80'h00_0060_00_0000_0C08_FFA4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2841_4 ( .OUT(na2841_2), .IN1(~na32_1), .IN2(na467_1), .IN3(na9180_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x75y75     80'h00_0060_00_0000_0C08_FFEA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2842_4 ( .OUT(na2842_2), .IN1(na155_1), .IN2(1'b0), .IN3(na354_2), .IN4(na9203_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y69     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2843_1 ( .OUT(na2843_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na88_1), .IN6(~na91_1), .IN7(~na90_1), .IN8(~na9162_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x66y95     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2844_4 ( .OUT(na2844_2), .IN1(na9699_2), .IN2(1'b1), .IN3(na2843_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x70y67     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2845_4 ( .OUT(na2845_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na797_1), .IN4(na2841_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y64     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2846_4 ( .OUT(na2846_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2843_1), .IN4(na2847_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x68y62     80'h00_0018_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2847_1 ( .OUT(na2847_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na155_1), .IN6(na2849_1), .IN7(1'b0), .IN8(na2841_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y73     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2848_4 ( .OUT(na2848_2), .IN1(na155_1), .IN2(~na2849_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x77y56     80'h00_0018_00_0040_0C6C_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2849_1 ( .OUT(na2849_1), .IN1(1'b0), .IN2(1'b1), .IN3(~na8096_2), .IN4(na5403_2), .IN5(~na356_2), .IN6(1'b1), .IN7(~na354_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y43     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2850_4 ( .OUT(na2850_2), .IN1(1'b1), .IN2(na2851_2), .IN3(na2843_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x71y64     80'h00_0060_00_0000_0C08_FFCD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2851_4 ( .OUT(na2851_2), .IN1(~na155_1), .IN2(na8097_2), .IN3(1'b0), .IN4(na2841_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x77y76     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2852_1 ( .OUT(na2852_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na155_1), .IN6(1'b0), .IN7(na8098_1), .IN8(na9337_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y45     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2853_1 ( .OUT(na2853_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2854_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2840_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y61     80'h00_0060_00_0000_0C08_FF12
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2854_4 ( .OUT(na2854_2), .IN1(na88_1), .IN2(~na91_1), .IN3(~na90_1), .IN4(~na9162_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y67     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2855_4 ( .OUT(na2855_2), .IN1(na2854_2), .IN2(1'b1), .IN3(na2845_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y64     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2856_1 ( .OUT(na2856_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2854_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2847_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x46y71     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2857_4 ( .OUT(na2857_2), .IN1(na2854_2), .IN2(na2851_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y73     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2858_1 ( .OUT(na2858_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na9698_2), .IN7(1'b1), .IN8(na2859_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x62y58     80'h00_0018_00_0000_0C88_41FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2859_1 ( .OUT(na2859_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na88_1), .IN6(~na91_1), .IN7(~na90_1), .IN8(na9162_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y75     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2860_4 ( .OUT(na2860_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2845_2), .IN4(na2859_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y36     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2861_1 ( .OUT(na2861_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9700_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2859_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y35     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2862_1 ( .OUT(na2862_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2851_2), .IN7(1'b1), .IN8(na2859_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y46     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2863_4 ( .OUT(na2863_2), .IN1(1'b1), .IN2(na2864_2), .IN3(1'b1), .IN4(na2840_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x57y62     80'h00_0060_00_0000_0C08_FF42
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2864_4 ( .OUT(na2864_2), .IN1(na88_1), .IN2(~na91_1), .IN3(~na90_1), .IN4(na9162_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y62     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2865_4 ( .OUT(na2865_2), .IN1(1'b1), .IN2(na2864_2), .IN3(na2845_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y63     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2866_1 ( .OUT(na2866_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2864_2), .IN7(1'b1), .IN8(na2847_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y79     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2867_4 ( .OUT(na2867_2), .IN1(1'b1), .IN2(na2864_2), .IN3(na9701_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y81     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2868_1 ( .OUT(na2868_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2869_1), .IN7(1'b1), .IN8(na2840_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x71y68     80'h00_0018_00_0000_0C88_21FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2869_1 ( .OUT(na2869_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na88_1), .IN6(~na91_1), .IN7(na90_1), .IN8(~na9162_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y74     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2870_4 ( .OUT(na2870_2), .IN1(1'b1), .IN2(na2869_1), .IN3(na2845_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y69     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2871_4 ( .OUT(na2871_2), .IN1(1'b1), .IN2(na2869_1), .IN3(1'b1), .IN4(na2847_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y63     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2872_1 ( .OUT(na2872_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2869_1), .IN7(na9701_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y54     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2873_1 ( .OUT(na2873_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2874_2), .IN8(na2840_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x84y57     80'h00_0060_00_0000_0C08_FF22
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2874_4 ( .OUT(na2874_2), .IN1(na88_1), .IN2(~na91_1), .IN3(na90_1), .IN4(~na9162_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2875_1 ( .OUT(na2875_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9699_2), .IN6(1'b1), .IN7(na2874_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y51     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2876_4 ( .OUT(na2876_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2874_2), .IN4(na2847_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y50     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2877_4 ( .OUT(na2877_2), .IN1(1'b1), .IN2(na2851_2), .IN3(na2874_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y50     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2878_4 ( .OUT(na2878_2), .IN1(1'b1), .IN2(na2879_1), .IN3(1'b1), .IN4(na2840_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x73y72     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2879_1 ( .OUT(na2879_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na88_1), .IN6(~na91_1), .IN7(na90_1), .IN8(na9162_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x58y92     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2880_4 ( .OUT(na2880_2), .IN1(1'b1), .IN2(na2879_1), .IN3(na2845_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y90     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2881_1 ( .OUT(na2881_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2879_1), .IN7(1'b1), .IN8(na2847_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y79     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2882_4 ( .OUT(na2882_2), .IN1(1'b1), .IN2(na2879_1), .IN3(na9701_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y66     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2883_1 ( .OUT(na2883_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2884_2), .IN7(1'b1), .IN8(na2840_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x77y70     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2884_4 ( .OUT(na2884_2), .IN1(na88_1), .IN2(~na91_1), .IN3(na90_1), .IN4(na9162_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y75     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2885_1 ( .OUT(na2885_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2884_2), .IN7(na2845_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y78     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2886_4 ( .OUT(na2886_2), .IN1(1'b1), .IN2(na2884_2), .IN3(1'b1), .IN4(na2847_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x70y83     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2887_1 ( .OUT(na2887_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2884_2), .IN7(na9701_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y57     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2888_4 ( .OUT(na2888_2), .IN1(1'b1), .IN2(na9698_2), .IN3(1'b1), .IN4(na2889_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y54     80'h00_0018_00_0000_0C88_14FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2889_1 ( .OUT(na2889_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na88_1), .IN6(na91_1), .IN7(~na90_1), .IN8(~na9162_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y38     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2890_1 ( .OUT(na2890_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2845_2), .IN8(na2889_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y36     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2891_4 ( .OUT(na2891_2), .IN1(na9700_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2889_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x54y55     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2892_4 ( .OUT(na2892_2), .IN1(1'b1), .IN2(na2851_2), .IN3(1'b1), .IN4(na2889_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x113y88     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2894_4 ( .OUT(na2894_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3546_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2894_5 ( .OUT(na2894_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2894_2_i) );
// C_MX4b/D///      x99y102     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2895_1 ( .OUT(na2895_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9704_2),
                      .IN8(na3751_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2895_2 ( .OUT(na2895_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2895_1_i) );
// C_AND*/D//AND*/D      x90y52     80'h00_FE00_80_0000_0387_5C3C
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2897_1 ( .OUT(na2897_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(~na4093_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2897_2 ( .OUT(na2897_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2897_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a2897_4 ( .OUT(na2897_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(1'b1), .IN4(~na4095_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a2897_5 ( .OUT(na2897_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2897_2_i) );
// C_AND/D//AND/D      x89y48     80'h00_FE00_80_0000_0C88_ACCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2898_1 ( .OUT(na2898_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(na4104_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2898_2 ( .OUT(na2898_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2898_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2898_4 ( .OUT(na2898_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(1'b1), .IN4(na4087_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2898_5 ( .OUT(na2898_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2898_2_i) );
// C_AND*/D//AND*/D      x88y47     80'h00_FE00_80_0000_0387_5C5C
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2899_1 ( .OUT(na2899_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(~na4104_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2899_2 ( .OUT(na2899_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2899_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a2899_4 ( .OUT(na2899_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(~na4093_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a2899_5 ( .OUT(na2899_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2899_2_i) );
// C_AND/D//AND/D      x91y47     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2900_1 ( .OUT(na2900_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(1'b1), .IN8(na4102_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2900_2 ( .OUT(na2900_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2900_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2900_4 ( .OUT(na2900_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(1'b1), .IN4(na4087_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2900_5 ( .OUT(na2900_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2900_2_i) );
// C_AND/D//AND/D      x88y50     80'h00_FE00_80_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2901_1 ( .OUT(na2901_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(1'b1), .IN8(na4102_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2901_2 ( .OUT(na2901_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2901_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2901_4 ( .OUT(na2901_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(na4100_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2901_5 ( .OUT(na2901_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2901_2_i) );
// C_AND*/D///      x89y51     80'h00_FE00_00_0000_0388_5CFF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a2902_1 ( .OUT(na2902_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(~na4100_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a2902_2 ( .OUT(na2902_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2902_1_i) );
// C_AND/D//AND/D      x87y50     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2904_1 ( .OUT(na2904_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(1'b1), .IN8(na4098_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2904_2 ( .OUT(na2904_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2904_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2904_4 ( .OUT(na2904_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(1'b1), .IN4(na4098_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2904_5 ( .OUT(na2904_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2904_2_i) );
// C_MX4b/D///      x119y87     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2906_1 ( .OUT(na2906_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2906_1), .IN6(na1099_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2906_2 ( .OUT(na2906_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2906_1_i) );
// C_AND/D//AND/D      x94y46     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2907_1 ( .OUT(na2907_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na172_2), .IN7(na4096_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2907_2 ( .OUT(na2907_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2907_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2907_4 ( .OUT(na2907_2_i), .IN1(1'b1), .IN2(na172_2), .IN3(na4096_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2907_5 ( .OUT(na2907_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2907_2_i) );
// C_MX4b/D///      x128y84     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2908_1 ( .OUT(na2908_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3056_1),
                      .IN8(na2908_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2908_2 ( .OUT(na2908_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2908_1_i) );
// C_MX4b/D///      x125y86     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2909_1 ( .OUT(na2909_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3058_1), .IN6(na2909_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2909_2 ( .OUT(na2909_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2909_1_i) );
// C_MX4b/D///      x119y86     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2910_1 ( .OUT(na2910_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9707_2), .IN6(na3060_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2910_2 ( .OUT(na2910_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2910_1_i) );
// C_MX4b/D///      x127y82     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2911_1 ( .OUT(na2911_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3062_1),
                      .IN8(na9708_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2911_2 ( .OUT(na2911_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2911_1_i) );
// C_MX4b/D///      x126y83     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2912_1 ( .OUT(na2912_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2912_1),
                      .IN8(na1445_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2912_2 ( .OUT(na2912_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2912_1_i) );
// C_MX4b/D///      x126y90     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2913_1 ( .OUT(na2913_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3068_1),
                      .IN8(na2913_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2913_2 ( .OUT(na2913_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2913_1_i) );
// C_MX4b/D///      x125y90     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2914_1 ( .OUT(na2914_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9711_2), .IN6(na3077_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2914_2 ( .OUT(na2914_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2914_1_i) );
// C_MX4b/D///      x127y88     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2915_1 ( .OUT(na2915_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9712_2),
                      .IN8(na3079_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2915_2 ( .OUT(na2915_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2915_1_i) );
// C_///AND/D      x89y47     80'h00_FE00_80_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2917_4 ( .OUT(na2917_2_i), .IN1(~na2917_2), .IN2(na172_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2917_5 ( .OUT(na2917_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2917_2_i) );
// C_AND/D///      x117y77     80'h00_FE00_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2918_1 ( .OUT(na2918_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10027_2), .IN6(~na9941_2), .IN7(na2932_1),
                      .IN8(na154_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2918_2 ( .OUT(na2918_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2918_1_i) );
// C_MX4b/D///      x121y102     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2919_1 ( .OUT(na2919_1_i), .IN1(na7054_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na8099_2), .IN6(na2919_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2919_2 ( .OUT(na2919_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2919_1_i) );
// C_///AND/D      x107y71     80'h00_FE00_80_0000_0C08_FF32
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2920_4 ( .OUT(na2920_2_i), .IN1(na8107_2), .IN2(~na2921_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2920_5 ( .OUT(na2920_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2920_2_i) );
// C_ORAND////      x107y72     80'h00_0018_00_0000_0C88_73FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2921_1 ( .OUT(na2921_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na6475_1), .IN7(~na2950_1), .IN8(~na2948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x121y64     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2922_1 ( .OUT(na2922_1_i), .IN1(~na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6484_1), .IN6(na2922_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2922_2 ( .OUT(na2922_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2922_1_i) );
// C_AND////      x113y79     80'h00_0018_00_0000_0C88_C1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2923_1 ( .OUT(na2923_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10027_2), .IN6(~na2931_1), .IN7(1'b1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x121y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2924_1 ( .OUT(na2924_1_i), .IN1(na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2924_1), .IN6(na6483_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2924_2 ( .OUT(na2924_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2924_1_i) );
// C_MX4b/D///      x121y67     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2925_1 ( .OUT(na2925_1_i), .IN1(na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2925_1), .IN6(na6482_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2925_2 ( .OUT(na2925_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2925_1_i) );
// C_MX4b/D///      x125y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2926_1 ( .OUT(na2926_1_i), .IN1(na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2926_1), .IN6(na6481_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2926_2 ( .OUT(na2926_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2926_1_i) );
// C_MX4b/D///      x121y68     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2927_1 ( .OUT(na2927_1_i), .IN1(~na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6480_1), .IN6(na2927_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2927_2 ( .OUT(na2927_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2927_1_i) );
// C_MX4b/D///      x127y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2928_1 ( .OUT(na2928_1_i), .IN1(na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2928_1), .IN6(na6479_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2928_2 ( .OUT(na2928_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2928_1_i) );
// C_MX4b/D///      x126y67     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2929_1 ( .OUT(na2929_1_i), .IN1(na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2929_1),
                      .IN8(na6478_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2929_2 ( .OUT(na2929_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2929_1_i) );
// C_MX4b/D///      x119y65     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2930_1 ( .OUT(na2930_1_i), .IN1(na2923_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2930_1), .IN6(na6477_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2930_2 ( .OUT(na2930_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2930_1_i) );
// C_AND/D///      x129y68     80'h00_FE00_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2931_1 ( .OUT(na2931_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2932_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2931_2 ( .OUT(na2931_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2931_1_i) );
// C_MX4a////      x114y83     80'h00_0018_00_0040_0C5C_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2932_1 ( .OUT(na2932_1), .IN1(1'b1), .IN2(1'b0), .IN3(~na8101_1), .IN4(na154_1), .IN5(1'b1), .IN6(na2931_1), .IN7(~na8101_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x123y100     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2933_4 ( .OUT(na2933_2_i), .IN1(na8103_1), .IN2(na2933_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2933_5 ( .OUT(na2933_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2933_2_i) );
// C_MX4b/D///      x87y90     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2935_1 ( .OUT(na2935_1_i), .IN1(~na212_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na8104_1), .IN6(na2935_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2935_2 ( .OUT(na2935_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2935_1_i) );
// C_MX4b/D///      x123y86     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2936_1 ( .OUT(na2936_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3081_1), .IN6(na2936_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2936_2 ( .OUT(na2936_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2936_1_i) );
// C_///ICOMP/D      x86y93     80'h00_FE00_80_0000_0C08_FF36
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2937_4 ( .OUT(na2937_2_i), .IN1(~na212_1), .IN2(na9715_2), .IN3(1'b0), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2937_5 ( .OUT(na2937_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2937_2_i) );
// C_MX4b/D///      x115y60     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2938_1 ( .OUT(na2938_1_i), .IN1(~na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6484_1), .IN6(na2938_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2938_2 ( .OUT(na2938_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2938_1_i) );
// C_MX4b/D///      x117y61     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2939_1 ( .OUT(na2939_1_i), .IN1(na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2939_1), .IN6(na6482_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2939_2 ( .OUT(na2939_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2939_1_i) );
// C_MX4b/D///      x119y59     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2940_1 ( .OUT(na2940_1_i), .IN1(na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2940_1), .IN6(na6481_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2940_2 ( .OUT(na2940_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2940_1_i) );
// C_MX4b/D///      x117y59     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2941_1 ( .OUT(na2941_1_i), .IN1(na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2941_1), .IN6(na6479_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2941_2 ( .OUT(na2941_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2941_1_i) );
// C_MX4b/D///      x120y57     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2942_1 ( .OUT(na2942_1_i), .IN1(na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2942_1),
                      .IN8(na6478_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2942_2 ( .OUT(na2942_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2942_1_i) );
// C_MX4b/D///      x126y86     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2943_1 ( .OUT(na2943_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3083_1),
                      .IN8(na2943_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2943_2 ( .OUT(na2943_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2943_1_i) );
// C_MX4b/D///      x125y88     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2944_1 ( .OUT(na2944_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9717_2), .IN6(na3085_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2944_2 ( .OUT(na2944_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2944_1_i) );
// C_MX4b/D///      x125y92     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2945_1 ( .OUT(na2945_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9718_2),
                      .IN8(na3087_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2945_2 ( .OUT(na2945_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2945_1_i) );
// C_MX4b/D///      x123y90     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2946_1 ( .OUT(na2946_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3089_1), .IN6(na2946_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2946_2 ( .OUT(na2946_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2946_1_i) );
// C_MX4b/D///      x113y59     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2947_1 ( .OUT(na2947_1_i), .IN1(na572_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2947_1), .IN6(na6477_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2947_2 ( .OUT(na2947_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2947_1_i) );
// C_///AND/D      x122y56     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2948_4 ( .OUT(na2948_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na2949_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2948_5 ( .OUT(na2948_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2948_2_i) );
// C_MX4a////      x114y67     80'h00_0018_00_0040_0CC9_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2949_1 ( .OUT(na2949_1), .IN1(na8107_2), .IN2(1'b0), .IN3(1'b1), .IN4(~na8106_1), .IN5(1'b1), .IN6(na2921_1), .IN7(1'b1),
                      .IN8(~na2948_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x120y53     80'h00_FE00_00_0040_0C0C_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2950_1 ( .OUT(na2950_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na2950_1), .IN4(na10028_2), .IN5(na8107_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na6626_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2950_2 ( .OUT(na2950_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2950_1_i) );
// C_///ORAND/D      x121y95     80'h00_FE00_80_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2951_4 ( .OUT(na2951_2_i), .IN1(na8109_2), .IN2(na2952_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2951_5 ( .OUT(na2951_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2951_2_i) );
// C_///AND/      x127y98     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2952_4 ( .OUT(na2952_2), .IN1(1'b1), .IN2(na3739_1), .IN3(1'b1), .IN4(~na654_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND/D      x126y96     80'h00_FE00_80_0000_0C88_3E3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2953_1 ( .OUT(na2953_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8111_2), .IN6(na2954_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2953_2 ( .OUT(na2953_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2953_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2953_4 ( .OUT(na2953_2_i), .IN1(na6935_1), .IN2(na657_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2953_5 ( .OUT(na2953_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2953_2_i) );
// C_///AND/      x125y98     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2954_4 ( .OUT(na2954_2), .IN1(na3737_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na654_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x125y76     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2955_1 ( .OUT(na2955_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9720_2), .IN6(na3091_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2955_2 ( .OUT(na2955_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2955_1_i) );
// C_MX4b/D///      x125y80     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2956_1 ( .OUT(na2956_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3093_1), .IN6(na2956_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2956_2 ( .OUT(na2956_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2956_1_i) );
// C_MX4b/D///      x123y78     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2957_1 ( .OUT(na2957_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9721_2),
                      .IN8(na3095_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2957_2 ( .OUT(na2957_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2957_1_i) );
// C_///AND/      x121y94     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2959_4 ( .OUT(na2959_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na9298_2), .IN4(~na753_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x91y89     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2960_1 ( .OUT(na2960_1_i), .IN1(1'b1), .IN2(na758_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2960_1), .IN6(na2961_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2960_2 ( .OUT(na2960_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2960_1_i) );
// C_AND////      x89y90     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2961_1 ( .OUT(na2961_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na7004_2), .IN6(1'b1), .IN7(na3871_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x99y68     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2962_1 ( .OUT(na2962_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na155_1), .IN6(na2962_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2962_2 ( .OUT(na2962_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2962_1_i) );
// C_MX4b/D///      x95y81     80'h00_FE00_00_0040_0A32_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2963_1 ( .OUT(na2963_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2963_1), .IN6(~na2852_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2963_2 ( .OUT(na2963_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2963_1_i) );
// C_MX4b/D///      x95y82     80'h00_FE00_00_0040_0A31_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2964_1 ( .OUT(na2964_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na2848_2), .IN6(na2964_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2964_2 ( .OUT(na2964_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2964_1_i) );
// C_MX4b/D///      x87y82     80'h00_FE00_00_0040_0A31_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2965_1 ( .OUT(na2965_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na2842_2), .IN6(na2965_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2965_2 ( .OUT(na2965_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2965_1_i) );
// C_MX4b/D///      x86y83     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2966_1 ( .OUT(na2966_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2551_2),
                      .IN8(na9722_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2966_2 ( .OUT(na2966_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2966_1_i) );
// C_MX4b/D///      x90y76     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2967_1 ( .OUT(na2967_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9723_2),
                      .IN8(na2549_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2967_2 ( .OUT(na2967_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2967_1_i) );
// C_MX4b/D///      x120y76     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2968_1 ( .OUT(na2968_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na2968_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2968_2 ( .OUT(na2968_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2968_1_i) );
// C_MX4b/D///      x87y70     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2969_1 ( .OUT(na2969_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2540_1), .IN6(na2969_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2969_2 ( .OUT(na2969_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2969_1_i) );
// C_MX4b/D///      x86y81     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2970_1 ( .OUT(na2970_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2970_1),
                      .IN8(na2528_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2970_2 ( .OUT(na2970_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2970_1_i) );
// C_MX4b/D///      x91y84     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2971_1 ( .OUT(na2971_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9724_2),
                      .IN8(na2526_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2971_2 ( .OUT(na2971_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2971_1_i) );
// C_AND/D//AND/D      x129y52     80'h00_FE00_80_0000_0C88_5553
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2972_1 ( .OUT(na2972_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2973_1), .IN6(1'b1), .IN7(~na986_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2972_2 ( .OUT(na2972_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2972_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2972_4 ( .OUT(na2972_2_i), .IN1(1'b1), .IN2(~na1108_1), .IN3(~na986_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2972_5 ( .OUT(na2972_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2972_2_i) );
// C_MX2b////      x129y49     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2973_1 ( .OUT(na2973_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na500_2), .IN5(1'b0), .IN6(~na2972_1), .IN7(1'b0), .IN8(~na8116_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x90y70     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2974_1 ( .OUT(na2974_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na5591_1), .IN6(na9727_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2974_2 ( .OUT(na2974_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2974_1_i) );
// C_MX4b/D///      x91y69     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2975_1 ( .OUT(na2975_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2975_1), .IN6(na5590_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2975_2 ( .OUT(na2975_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2975_1_i) );
// C_MX4b/D///      x88y78     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2976_1 ( .OUT(na2976_1_i), .IN1(na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na5589_1),
                      .IN8(na2976_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2976_2 ( .OUT(na2976_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2976_1_i) );
// C_MX4b/D///      x93y73     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2977_1 ( .OUT(na2977_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2977_1), .IN6(na5588_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2977_2 ( .OUT(na2977_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2977_1_i) );
// C_MX4b/D///      x88y81     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2978_1 ( .OUT(na2978_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na2978_1),
                      .IN8(na5587_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2978_2 ( .OUT(na2978_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2978_1_i) );
// C_MX4b/D///      x88y72     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2979_1 ( .OUT(na2979_1_i), .IN1(~na421_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9729_2), .IN6(na5586_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2979_2 ( .OUT(na2979_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2979_1_i) );
// C_///AND/D      x104y70     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2980_4 ( .OUT(na2980_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1132_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a2980_5 ( .OUT(na2980_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2980_2_i) );
// C_ORAND/D///      x121y69     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2981_1 ( .OUT(na2981_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8118_1), .IN6(na2982_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2981_2 ( .OUT(na2981_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2981_1_i) );
// C_///AND/      x127y68     80'h00_0060_00_0000_0C08_FF24
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2982_4 ( .OUT(na2982_2), .IN1(~na155_1), .IN2(na647_1), .IN3(na224_1), .IN4(~na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x115y94     80'h00_FE00_00_0040_0C0A_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2983_1 ( .OUT(na2983_1_i), .IN1(1'b0), .IN2(na2983_1), .IN3(1'b0), .IN4(na8119_2), .IN5(~na9940_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na2984_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2983_2 ( .OUT(na2983_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2983_1_i) );
// C_ORAND////      x116y98     80'h00_0018_00_0000_0888_F575
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2984_1 ( .OUT(na2984_1), .IN1(~na951_1), .IN2(1'b0), .IN3(~na2986_1), .IN4(~na8121_1), .IN5(~na951_2), .IN6(1'b0), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x112y105     80'h00_FE18_00_0000_0666_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2986_1 ( .OUT(na2986_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2987_1), .IN6(~na2983_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2986_5 ( .OUT(na2986_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2986_1) );
// C_MX4b/D///      x115y97     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2987_1 ( .OUT(na2987_1_i), .IN1(1'b1), .IN2(~na2983_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2987_1), .IN6(na8123_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2987_2 ( .OUT(na2987_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2987_1_i) );
// C_ORAND/D///      x100y88     80'h00_FE00_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2989_1 ( .OUT(na2989_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8125_2), .IN6(na2990_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2989_2 ( .OUT(na2989_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2989_1_i) );
// C_///ORAND/      x93y94     80'h00_0060_00_0000_0C08_FFC7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2990_4 ( .OUT(na2990_2), .IN1(~na1225_1), .IN2(~na1173_1), .IN3(1'b0), .IN4(na2989_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x105y61     80'h00_FE00_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2991_1 ( .OUT(na2991_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9414_2), .IN6(~na7097_1), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2991_2 ( .OUT(na2991_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2991_1_i) );
// C_MX4b/D///      x101y61     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2992_1 ( .OUT(na2992_1_i), .IN1(1'b1), .IN2(na1130_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2992_1), .IN6(na3841_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2992_2 ( .OUT(na2992_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2992_1_i) );
// C_MX4b/D///      x103y62     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2993_1 ( .OUT(na2993_1_i), .IN1(1'b1), .IN2(~na1130_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3839_2), .IN6(na2993_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2993_2 ( .OUT(na2993_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2993_1_i) );
// C_MX4b/D///      x85y83     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2994_1 ( .OUT(na2994_1_i), .IN1(na2680_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2994_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2994_2 ( .OUT(na2994_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2994_1_i) );
// C_MX4b/D///      x104y61     80'h00_FE00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2995_1 ( .OUT(na2995_1_i), .IN1(1'b1), .IN2(~na1130_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3839_1), .IN6(na9731_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2995_2 ( .OUT(na2995_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2995_1_i) );
// C_MX4b/D///      x99y63     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2996_1 ( .OUT(na2996_1_i), .IN1(1'b1), .IN2(na1130_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na2996_1), .IN6(~na9732_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a2996_2 ( .OUT(na2996_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2996_1_i) );
// C_MX4a////      x107y52     80'h00_0018_00_0040_0CF6_5300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2998_1 ( .OUT(na2998_1), .IN1(1'b1), .IN2(~na4108_1), .IN3(~na3849_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1130_1), .IN7(~na1136_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x109y50     80'h00_0018_00_0040_0CF9_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3000_1 ( .OUT(na3000_1), .IN1(~na4106_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na3847_2), .IN5(1'b1), .IN6(na1130_1), .IN7(~na1136_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x123y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3001_1 ( .OUT(na3001_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3001_1), .IN6(na1211_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3001_2 ( .OUT(na3001_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3001_1_i) );
// C_AND/D///      x50y109     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3002_1 ( .OUT(na3002_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3816_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3002_2 ( .OUT(na3002_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3002_1_i) );
// C_AND*/D//AND*/D      x123y45     80'h00_FE00_80_0000_0387_C3C3
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a3003_1 ( .OUT(na3003_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3778_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3003_2 ( .OUT(na3003_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3003_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a3003_4 ( .OUT(na3003_2_i), .IN1(1'b1), .IN2(~na3778_1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3003_5 ( .OUT(na3003_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3003_2_i) );
// C_AND*/D//AND/D      x125y43     80'h00_FE00_80_0000_0388_C3CC
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a3006_1 ( .OUT(na3006_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3774_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3006_2 ( .OUT(na3006_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3006_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3006_4 ( .OUT(na3006_2_i), .IN1(1'b1), .IN2(na3774_1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3006_5 ( .OUT(na3006_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3006_2_i) );
// C_MX4b/D///      x126y78     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3008_1 ( .OUT(na3008_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3097_1),
                      .IN8(na3008_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3008_2 ( .OUT(na3008_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3008_1_i) );
// C_MX4b/D///      x127y78     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3009_1 ( .OUT(na3009_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3099_1), .IN6(na3009_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3009_2 ( .OUT(na3009_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3009_1_i) );
// C_MX4b/D///      x123y76     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3010_1 ( .OUT(na3010_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9734_2),
                      .IN8(na3101_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3010_2 ( .OUT(na3010_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3010_1_i) );
// C_MX4b/D///      x121y78     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3011_1 ( .OUT(na3011_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3103_1),
                      .IN8(na9735_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3011_2 ( .OUT(na3011_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3011_1_i) );
// C_MX4b/D///      x123y77     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3012_1 ( .OUT(na3012_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3012_1), .IN6(na3105_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3012_2 ( .OUT(na3012_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3012_1_i) );
// C_///AND/D      x129y75     80'h00_FE00_80_0000_0C08_FF38
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3013_4 ( .OUT(na3013_2_i), .IN1(na9361_2), .IN2(na459_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3013_5 ( .OUT(na3013_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3013_2_i) );
// C_///AND/D      x102y79     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3014_4 ( .OUT(na3014_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3015_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3014_5 ( .OUT(na3014_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3014_2_i) );
// C_MX2a////      x112y75     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3015_1 ( .OUT(na3015_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na3014_2), .IN4(~na159_1), .IN5(na9235_2), .IN6(na955_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x106y78     80'h00_FE00_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3016_1 ( .OUT(na3016_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na906_1), .IN6(na459_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3016_2 ( .OUT(na3016_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3016_1_i) );
// C_MX4b/D///      x122y94     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3017_1 ( .OUT(na3017_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9736_2), .IN6(na1211_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3017_2 ( .OUT(na3017_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3017_1_i) );
// C_AND*/D//AND*/D      x126y43     80'h00_FE00_80_0000_0387_C5C5
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a3018_1 ( .OUT(na3018_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3804_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3018_2 ( .OUT(na3018_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3018_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a3018_4 ( .OUT(na3018_2_i), .IN1(~na3804_1), .IN2(1'b1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3018_5 ( .OUT(na3018_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3018_2_i) );
// C_AND*/D//AND*/D      x125y42     80'h00_FE00_80_0000_0387_C3C3
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a3020_1 ( .OUT(na3020_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3802_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3020_2 ( .OUT(na3020_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3020_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a3020_4 ( .OUT(na3020_2_i), .IN1(1'b1), .IN2(~na3802_1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3020_5 ( .OUT(na3020_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3020_2_i) );
// C_AND*/D//AND*/D      x126y42     80'h00_FE00_80_0000_0387_C5C5
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a3022_1 ( .OUT(na3022_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3800_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3022_2 ( .OUT(na3022_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3022_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a3022_4 ( .OUT(na3022_2_i), .IN1(~na3800_1), .IN2(1'b1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3022_5 ( .OUT(na3022_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3022_2_i) );
// C_AND/D//AND*/D      x124y41     80'h00_FE00_80_0000_0C87_CCC3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3024_1 ( .OUT(na3024_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3798_2), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3024_2 ( .OUT(na3024_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3024_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a3024_4 ( .OUT(na3024_2_i), .IN1(1'b1), .IN2(~na3798_1), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3024_5 ( .OUT(na3024_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3024_2_i) );
// C_AND/D//AND*/D      x123y42     80'h00_FE00_80_0000_0C87_CACC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3026_1 ( .OUT(na3026_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3783_2), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3026_2 ( .OUT(na3026_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3026_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a3026_4 ( .OUT(na3026_2_i), .IN1(1'b1), .IN2(na3026_2), .IN3(1'b1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3026_5 ( .OUT(na3026_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3026_2_i) );
// C_AND/D///      x126y40     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3027_1 ( .OUT(na3027_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3783_1), .IN6(1'b1), .IN7(1'b1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3027_2 ( .OUT(na3027_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3027_1_i) );
// C_///AND/D      x115y80     80'h00_FE00_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3029_4 ( .OUT(na3029_2_i), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3029_5 ( .OUT(na3029_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3029_2_i) );
// C_AND/D//AND/D      x119y50     80'h00_F600_80_0000_0C88_8C8A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3031_1 ( .OUT(na3031_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4075_2), .IN7(na1223_1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3031_2 ( .OUT(na3031_1), .CLK(na4116_1), .EN(~na57_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3031_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3031_4 ( .OUT(na3031_2_i), .IN1(na4077_1), .IN2(1'b1), .IN3(na1223_1), .IN4(na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3031_5 ( .OUT(na3031_2), .CLK(na4116_1), .EN(~na57_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3031_2_i) );
// C_AND/D//AND/D      x120y50     80'h00_F600_80_0000_0C88_8C2C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3032_1 ( .OUT(na3032_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4075_1), .IN7(na1223_1), .IN8(na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3032_2 ( .OUT(na3032_1), .CLK(na4116_1), .EN(~na57_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3032_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3032_4 ( .OUT(na3032_2_i), .IN1(1'b1), .IN2(na9365_2), .IN3(na1223_1), .IN4(~na3032_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3032_5 ( .OUT(na3032_2), .CLK(na4116_1), .EN(~na57_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3032_2_i) );
// C_MX4b/D///      x113y87     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3034_1 ( .OUT(na3034_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3001_1), .IN6(~na3035_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3034_2 ( .OUT(na3034_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3034_1_i) );
// C_MX2b////      x127y86     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3035_1 ( .OUT(na3035_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9737_2), .IN8(~na4055_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x114y89     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3036_1 ( .OUT(na3036_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2239_1), .IN6(~na3037_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3036_2 ( .OUT(na3036_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3036_1_i) );
// C_MX2b////      x119y94     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3037_1 ( .OUT(na3037_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4052_2), .IN8(~na3070_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x113y92     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3038_1 ( .OUT(na3038_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na990_1), .IN6(~na3039_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3038_2 ( .OUT(na3038_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3038_1_i) );
// C_MX2b////      x119y90     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3039_1 ( .OUT(na3039_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4052_1), .IN8(~na3071_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x117y87     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3040_1 ( .OUT(na3040_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1883_1), .IN6(~na3041_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3040_2 ( .OUT(na3040_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3040_1_i) );
// C_MX2b////      x117y90     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3041_1 ( .OUT(na3041_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9743_2), .IN8(~na4050_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x116y91     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3042_1 ( .OUT(na3042_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1868_1), .IN6(~na3043_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3042_2 ( .OUT(na3042_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3042_1_i) );
// C_MX2b////      x117y92     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3043_1 ( .OUT(na3043_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9745_2), .IN8(~na4050_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x117y85     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3044_1 ( .OUT(na3044_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1138_1), .IN6(~na3045_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3044_2 ( .OUT(na3044_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3044_1_i) );
// C_MX2b////      x119y92     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3045_1 ( .OUT(na3045_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4048_2), .IN8(~na3074_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x115y82     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3046_1 ( .OUT(na3046_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1869_1), .IN6(~na3047_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3046_2 ( .OUT(na3046_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3046_1_i) );
// C_MX2b////      x121y92     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3047_1 ( .OUT(na3047_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4048_1), .IN8(~na3075_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x114y92     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3048_1 ( .OUT(na3048_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2906_1), .IN6(~na3049_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3048_2 ( .OUT(na3048_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3048_1_i) );
// C_MX2b////      x121y76     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3049_1 ( .OUT(na3049_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9749_2), .IN8(~na4046_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x127y90     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3050_1 ( .OUT(na3050_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3212_1), .IN6(~na3051_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3050_2 ( .OUT(na3050_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3050_1_i) );
// C_MX2b////      x117y82     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3051_1 ( .OUT(na3051_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3116_1), .IN8(~na4046_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x128y86     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3052_1 ( .OUT(na3052_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2246_1), .IN6(~na3053_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3052_2 ( .OUT(na3052_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3052_1_i) );
// C_MX2b////      x117y88     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3053_1 ( .OUT(na3053_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4044_2), .IN8(~na3117_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x128y90     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3054_1 ( .OUT(na3054_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2254_1), .IN6(~na3055_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3054_2 ( .OUT(na3054_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3054_1_i) );
// C_MX2b////      x121y82     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3055_1 ( .OUT(na3055_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4044_1), .IN8(~na3123_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x116y81     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3056_1 ( .OUT(na3056_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2717_1), .IN6(~na3057_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3056_2 ( .OUT(na3056_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3056_1_i) );
// C_MX2a////      x125y84     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3057_1 ( .OUT(na3057_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na3124_1), .IN4(~na4041_2), .IN5(1'b1), .IN6(~na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x115y81     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3058_1 ( .OUT(na3058_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2745_1), .IN6(~na3059_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3058_2 ( .OUT(na3058_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3058_1_i) );
// C_MX2a////      x121y84     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3059_1 ( .OUT(na3059_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na3128_1), .IN4(~na4041_1), .IN5(1'b1), .IN6(~na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x117y94     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3060_1 ( .OUT(na3060_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na471_1), .IN6(~na3061_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3060_2 ( .OUT(na3060_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3060_1_i) );
// C_MX2a////      x117y84     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3061_1 ( .OUT(na3061_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4039_2), .IN4(~na3129_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x118y81     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3062_1 ( .OUT(na3062_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1726_1), .IN6(~na3063_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3062_2 ( .OUT(na3062_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3062_1_i) );
// C_MX2a////      x123y96     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3063_1 ( .OUT(na3063_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4039_1), .IN4(~na579_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x51y112     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3064_1 ( .OUT(na3064_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3835_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3064_2 ( .OUT(na3064_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3064_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3064_4 ( .OUT(na3064_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3835_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3064_5 ( .OUT(na3064_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3064_2_i) );
// C_MX4b/D///      x111y56     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3065_1 ( .OUT(na3065_1_i), .IN1(~na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6484_1), .IN6(na3065_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3065_2 ( .OUT(na3065_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3065_1_i) );
// C_MX4b/D///      x120y78     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3066_1 ( .OUT(na3066_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na261_1),
                      .IN8(na3066_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3066_2 ( .OUT(na3066_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3066_1_i) );
// C_MX4b/D///      x128y95     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3068_1 ( .OUT(na3068_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3211_1), .IN6(~na3069_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3068_2 ( .OUT(na3068_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3068_1_i) );
// C_MX2a////      x119y82     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3069_1 ( .OUT(na3069_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na791_1), .IN4(~na4037_1), .IN5(1'b1), .IN6(~na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x114y96     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3070_1 ( .OUT(na3070_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9740_2), .IN6(na1110_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3070_2 ( .OUT(na3070_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3070_1_i) );
// C_MX4b/D///      x118y96     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3071_1 ( .OUT(na3071_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9741_2), .IN6(na991_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3071_2 ( .OUT(na3071_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3071_1_i) );
// C_MX4b/D///      x114y88     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3072_1 ( .OUT(na3072_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9742_2), .IN6(na1105_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3072_2 ( .OUT(na3072_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3072_1_i) );
// C_MX4b/D///      x116y94     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3073_1 ( .OUT(na3073_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9744_2), .IN6(na1103_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3073_2 ( .OUT(na3073_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3073_1_i) );
// C_MX4b/D///      x118y94     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3074_1 ( .OUT(na3074_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1139_1), .IN6(na9746_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3074_2 ( .OUT(na3074_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3074_1_i) );
// C_MX4b/D///      x114y90     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3075_1 ( .OUT(na3075_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9747_2), .IN6(na1101_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3075_2 ( .OUT(na3075_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3075_1_i) );
// C_MX4b/D///      x116y90     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3076_1 ( .OUT(na3076_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9748_2), .IN6(na1099_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3076_2 ( .OUT(na3076_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3076_1_i) );
// C_MX4b/D///      x125y94     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3077_1 ( .OUT(na3077_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3203_1), .IN6(~na3078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3077_2 ( .OUT(na3077_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3077_1_i) );
// C_MX2a////      x127y92     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3078_1 ( .OUT(na3078_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4035_2), .IN4(~na832_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x128y92     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3079_1 ( .OUT(na3079_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3196_1), .IN6(~na3080_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3079_2 ( .OUT(na3079_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3079_1_i) );
// C_MX2a////      x119y88     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3080_1 ( .OUT(na3080_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4035_1), .IN4(~na1382_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x127y91     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3081_1 ( .OUT(na3081_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3193_1), .IN6(~na3082_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3081_2 ( .OUT(na3081_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3081_1_i) );
// C_MX2b////      x123y88     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3082_1 ( .OUT(na3082_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9517_2), .IN8(~na4033_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x126y89     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3083_1 ( .OUT(na3083_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3171_1), .IN6(~na3084_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3083_2 ( .OUT(na3083_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3083_1_i) );
// C_MX2a////      x123y84     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3084_1 ( .OUT(na3084_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2762_1), .IN4(~na4033_1), .IN5(1'b1), .IN6(~na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x117y80     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3085_1 ( .OUT(na3085_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3166_1), .IN6(~na3086_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3085_2 ( .OUT(na3085_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3085_1_i) );
// C_MX2a////      x115y78     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3086_1 ( .OUT(na3086_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4062_2), .IN4(~na2661_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x114y80     80'h00_FE00_00_0040_0A31_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3087_1 ( .OUT(na3087_1_i), .IN1(1'b1), .IN2(~na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(~na3088_1), .IN6(na3152_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3087_2 ( .OUT(na3087_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3087_1_i) );
// C_MX2a////      x123y93     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3088_1 ( .OUT(na3088_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4062_1), .IN4(~na3189_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x129y95     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3089_1 ( .OUT(na3089_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3150_1), .IN6(~na3090_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3089_2 ( .OUT(na3089_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3089_1_i) );
// C_MX2a////      x133y90     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3090_1 ( .OUT(na3090_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na3183_1), .IN4(~na4060_2), .IN5(1'b1), .IN6(~na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x127y80     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3091_1 ( .OUT(na3091_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na2156_1), .IN6(~na3092_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3091_2 ( .OUT(na3091_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3091_1_i) );
// C_MX2b////      x131y84     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3092_1 ( .OUT(na3092_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9780_2), .IN8(~na4060_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x129y79     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3093_1 ( .OUT(na3093_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1889_1), .IN6(~na3094_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3093_2 ( .OUT(na3093_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3093_1_i) );
// C_MX2b////      x131y82     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3094_1 ( .OUT(na3094_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4058_2), .IN8(~na3165_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x132y80     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3095_1 ( .OUT(na3095_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3136_1), .IN6(~na3096_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3095_2 ( .OUT(na3095_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3095_1_i) );
// C_MX2b////      x133y80     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3096_1 ( .OUT(na3096_1), .IN1(1'b1), .IN2(na1447_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4058_1), .IN8(~na3156_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x114y79     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3097_1 ( .OUT(na3097_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1697_1), .IN6(~na3098_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3097_2 ( .OUT(na3097_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3097_1_i) );
// C_MX2a////      x123y82     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3098_1 ( .OUT(na3098_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na3155_1), .IN4(~na4056_2), .IN5(1'b1), .IN6(~na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x127y79     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3099_1 ( .OUT(na3099_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na1658_1), .IN6(~na3100_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3099_2 ( .OUT(na3099_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3099_1_i) );
// C_MX2a////      x121y80     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3100_1 ( .OUT(na3100_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na9739_2), .IN4(~na4056_1), .IN5(1'b1), .IN6(~na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x130y78     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3101_1 ( .OUT(na3101_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3121_1), .IN6(~na3102_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3101_2 ( .OUT(na3101_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3101_1_i) );
// C_MX2a////      x119y80     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3102_1 ( .OUT(na3102_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4042_2), .IN4(~na2968_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x128y77     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3103_1 ( .OUT(na3103_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(na6626_1), .IN5(na3114_1), .IN6(~na3104_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3103_2 ( .OUT(na3103_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3103_1_i) );
// C_MX2a////      x121y90     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3104_1 ( .OUT(na3104_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na4042_1), .IN4(~na2168_1), .IN5(1'b1), .IN6(na1447_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x129y78     80'h00_FE00_00_0040_0AC8_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3105_1 ( .OUT(na3105_1_i), .IN1(1'b1), .IN2(na3178_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1892_1),
                      .IN8(~na3106_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3105_2 ( .OUT(na3105_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3105_1_i) );
// C_MX2b////      x124y80     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3106_1 ( .OUT(na3106_1), .IN1(1'b1), .IN2(~na1447_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na9538_2), .IN6(na3105_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//AND/D      x87y84     80'h00_FE00_80_0000_0C88_3E8F
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3107_1 ( .OUT(na3107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8134_2), .IN6(na3108_2), .IN7(1'b0), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3107_2 ( .OUT(na3107_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3107_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3107_4 ( .OUT(na3107_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3186_2), .IN4(na9750_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3107_5 ( .OUT(na3107_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3107_2_i) );
// C_///ORAND/      x99y96     80'h00_0060_00_0000_0C08_FF7C
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3108_4 ( .OUT(na3108_2), .IN1(1'b0), .IN2(na3107_1), .IN3(~na1312_1), .IN4(~na3016_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x121y88     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3109_1 ( .OUT(na3109_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3034_1), .IN6(na3109_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3109_2 ( .OUT(na3109_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3109_1_i) );
// C_MX4b/D///      x123y94     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3110_1 ( .OUT(na3110_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3036_1),
                      .IN8(na9752_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3110_2 ( .OUT(na3110_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3110_1_i) );
// C_MX4b/D///      x123y92     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3111_1 ( .OUT(na3111_1_i), .IN1(na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9753_2), .IN6(na3038_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3111_2 ( .OUT(na3111_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3111_1_i) );
// C_MX4b/D///      x121y86     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3112_1 ( .OUT(na3112_1_i), .IN1(~na3013_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3040_1), .IN6(na3112_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3112_2 ( .OUT(na3112_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3112_1_i) );
// C_MX4b/D///      x100y99     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3113_1 ( .OUT(na3113_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3113_1),
                      .IN8(na3744_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3113_2 ( .OUT(na3113_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3113_1_i) );
// C_MX4b/D///      x115y75     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3114_1 ( .OUT(na3114_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3114_1), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3114_2 ( .OUT(na3114_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3114_1_i) );
// C_AND/D//AND/D      x52y116     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3115_1 ( .OUT(na3115_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3815_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3115_2 ( .OUT(na3115_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3115_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3115_4 ( .OUT(na3115_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3815_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3115_5 ( .OUT(na3115_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3115_2_i) );
// C_MX4b/D///      x120y87     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3116_1 ( .OUT(na3116_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3116_1),
                      .IN8(na1097_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3116_2 ( .OUT(na3116_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3116_1_i) );
// C_MX4b/D///      x120y86     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3117_1 ( .OUT(na3117_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1095_2),
                      .IN8(na3117_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3117_2 ( .OUT(na3117_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3117_1_i) );
// C_MX4b/D///      x91y97     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3118_1 ( .OUT(na3118_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9755_2),
                      .IN8(na3744_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3118_2 ( .OUT(na3118_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3118_1_i) );
// C_MX4b/D///      x100y100     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3119_1 ( .OUT(na3119_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3746_1),
                      .IN8(na3119_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3119_2 ( .OUT(na3119_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3119_1_i) );
// C_MX4b/D///      x119y71     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3121_1 ( .OUT(na3121_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na9756_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3121_2 ( .OUT(na3121_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3121_1_i) );
// C_AND/D//AND/D      x50y116     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3122_1 ( .OUT(na3122_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3818_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3122_2 ( .OUT(na3122_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3122_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3122_4 ( .OUT(na3122_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(na3818_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3122_5 ( .OUT(na3122_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3122_2_i) );
// C_MX4b/D///      x120y90     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3123_1 ( .OUT(na3123_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9757_2), .IN6(na993_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3123_2 ( .OUT(na3123_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3123_1_i) );
// C_MX4b/D///      x120y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3124_1 ( .OUT(na3124_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9758_2), .IN6(na961_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3124_2 ( .OUT(na3124_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3124_1_i) );
// C_MX4b/D///      x119y64     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3125_1 ( .OUT(na3125_1_i), .IN1(~na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6484_1), .IN6(na3125_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3125_2 ( .OUT(na3125_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3125_1_i) );
// C_MX4b/D///      x101y108     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3126_1 ( .OUT(na3126_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3746_2),
                      .IN8(na9760_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3126_2 ( .OUT(na3126_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3126_1_i) );
// C_AND/D//AND/D      x50y117     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3127_1 ( .OUT(na3127_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3820_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3127_2 ( .OUT(na3127_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3127_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3127_4 ( .OUT(na3127_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3820_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3127_5 ( .OUT(na3127_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3127_2_i) );
// C_MX4b/D///      x118y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3128_1 ( .OUT(na3128_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9761_2), .IN6(na1091_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3128_2 ( .OUT(na3128_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3128_1_i) );
// C_MX4b/D///      x118y92     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3129_1 ( .OUT(na3129_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9763_2), .IN6(na472_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3129_2 ( .OUT(na3129_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3129_1_i) );
// C_MX4b/D///      x96y96     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3130_1 ( .OUT(na3130_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3742_1),
                      .IN8(na3130_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3130_2 ( .OUT(na3130_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3130_1_i) );
// C_AND/D//AND/D      x52y118     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3131_1 ( .OUT(na3131_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3822_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3131_2 ( .OUT(na3131_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3131_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3131_4 ( .OUT(na3131_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(na3822_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3131_5 ( .OUT(na3131_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3131_2_i) );
// C_MX4b/D///      x113y91     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3132_1 ( .OUT(na3132_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3132_1), .IN6(na1105_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a3132_2 ( .OUT(na3132_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3132_1_i) );
// C_MX4b/D///      x104y107     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3134_1 ( .OUT(na3134_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3134_1),
                      .IN8(na3748_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3134_2 ( .OUT(na3134_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3134_1_i) );
// C_MX4b/D///      x117y81     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3136_1 ( .OUT(na3136_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na9765_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3136_2 ( .OUT(na3136_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3136_1_i) );
// C_AND/D//AND/D      x49y117     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3137_1 ( .OUT(na3137_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3824_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3137_2 ( .OUT(na3137_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3137_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3137_4 ( .OUT(na3137_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3824_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3137_5 ( .OUT(na3137_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3137_2_i) );
// C_MX4b/D///      x91y96     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3138_1 ( .OUT(na3138_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9766_2),
                      .IN8(na3771_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3138_2 ( .OUT(na3138_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3138_1_i) );
// C_MX4b/D///      x106y106     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3139_1 ( .OUT(na3139_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3750_1),
                      .IN8(na3139_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3139_2 ( .OUT(na3139_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3139_1_i) );
// C_AND/D///      x106y71     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3140_1 ( .OUT(na3140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na9359_2), .IN7(1'b1), .IN8(na949_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3140_2 ( .OUT(na3140_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3140_1_i) );
// C_MX4b/D///      x100y97     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3141_1 ( .OUT(na3141_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3769_2),
                      .IN8(na9767_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3141_2 ( .OUT(na3141_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3141_1_i) );
// C_///AND*/D      x51y119     80'h00_FE00_80_0000_0C07_FF3A
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a3142_4 ( .OUT(na3142_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3829_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3142_5 ( .OUT(na3142_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3142_2_i) );
// C_AND/D///      x84y84     80'h00_FE00_00_0000_0888_C8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3143_1 ( .OUT(na3143_1_i), .IN1(na4855_2), .IN2(na435_2), .IN3(1'b1), .IN4(1'b1), .IN5(na9954_2), .IN6(na435_1), .IN7(1'b1),
                      .IN8(na9223_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3143_2 ( .OUT(na3143_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3143_1_i) );
// C_AND/D///      x90y88     80'h00_FE00_00_0000_0888_F8A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3145_1 ( .OUT(na3145_1_i), .IN1(na428_1), .IN2(na435_1), .IN3(na433_1), .IN4(1'b1), .IN5(na9954_2), .IN6(na927_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3145_2 ( .OUT(na3145_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3145_1_i) );
// C_MX4b/D///      x92y96     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3146_1 ( .OUT(na3146_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3769_1),
                      .IN8(na3146_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3146_2 ( .OUT(na3146_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3146_1_i) );
// C_MX4b/D///      x100y107     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3147_1 ( .OUT(na3147_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3147_1),
                      .IN8(na3753_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3147_2 ( .OUT(na3147_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3147_1_i) );
// C_MX4b/D///      x95y96     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3148_1 ( .OUT(na3148_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9768_2),
                      .IN8(na3767_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3148_2 ( .OUT(na3148_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3148_1_i) );
// C_AND/D///      x88y89     80'h00_FE00_00_0000_0888_A2F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3149_1 ( .OUT(na3149_1_i), .IN1(na428_2), .IN2(na1880_2), .IN3(1'b1), .IN4(1'b1), .IN5(na428_1), .IN6(~na435_1), .IN7(na433_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3149_2 ( .OUT(na3149_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3149_1_i) );
// C_MX4b/D///      x115y95     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3150_1 ( .OUT(na3150_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3150_1), .IN6(na1073_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3150_2 ( .OUT(na3150_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3150_1_i) );
// C_MX4b/D///      x98y100     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3151_1 ( .OUT(na3151_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9769_2),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3151_2 ( .OUT(na3151_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3151_1_i) );
// C_MX4b/D///      x115y102     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3152_1 ( .OUT(na3152_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na3152_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3152_2 ( .OUT(na3152_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3152_1_i) );
// C_MX4b/D///      x106y98     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3153_1 ( .OUT(na3153_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9771_2), .IN6(na259_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3153_2 ( .OUT(na3153_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3153_1_i) );
// C_MX4b/D///      x112y56     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3154_1 ( .OUT(na3154_1_i), .IN1(na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9772_2), .IN6(na6483_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3154_2 ( .OUT(na3154_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3154_1_i) );
// C_MX4b/D///      x118y79     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3155_1 ( .OUT(na3155_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9773_2), .IN6(na262_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3155_2 ( .OUT(na3155_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3155_1_i) );
// C_MX4b/D///      x120y82     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3156_1 ( .OUT(na3156_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1),
                      .IN8(na3156_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3156_2 ( .OUT(na3156_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3156_1_i) );
// C_MX4b/D///      x103y103     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3158_1 ( .OUT(na3158_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3158_1), .IN6(na991_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3158_2 ( .OUT(na3158_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3158_1_i) );
// C_AND/D//AND/D      x49y111     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3159_1 ( .OUT(na3159_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3837_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3159_2 ( .OUT(na3159_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3159_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3159_4 ( .OUT(na3159_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(na3837_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3159_5 ( .OUT(na3159_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3159_2_i) );
// C_MX4b/D///      x103y105     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3161_1 ( .OUT(na3161_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3161_1), .IN6(na1110_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3161_2 ( .OUT(na3161_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3161_1_i) );
// C_AND/D//AND/D      x50y113     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3162_1 ( .OUT(na3162_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3807_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3162_2 ( .OUT(na3162_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3162_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3162_4 ( .OUT(na3162_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3807_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3162_5 ( .OUT(na3162_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3162_2_i) );
// C_MX4b/D///      x112y58     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3163_1 ( .OUT(na3163_1_i), .IN1(na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9775_2), .IN6(na6482_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3163_2 ( .OUT(na3163_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3163_1_i) );
// C_MX4b/D///      x114y58     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3164_1 ( .OUT(na3164_1_i), .IN1(na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9776_2), .IN6(na6481_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3164_2 ( .OUT(na3164_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3164_1_i) );
// C_MX4b/D///      x118y84     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3165_1 ( .OUT(na3165_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na264_1),
                      .IN8(na3165_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3165_2 ( .OUT(na3165_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3165_1_i) );
// C_MX4b/D///      x117y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3166_1 ( .OUT(na3166_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3166_1), .IN6(na454_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3166_2 ( .OUT(na3166_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3166_1_i) );
// C_AND/D///      x105y100     80'h00_F900_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3167_1 ( .OUT(na3167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na6065_2), .IN7(na933_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3167_2 ( .OUT(na3167_1), .CLK(~na4116_1), .EN(na3237_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3167_1_i) );
// C_MX4b/D///      x108y88     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3168_1 ( .OUT(na3168_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na260_1),
                      .IN8(na3168_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3168_2 ( .OUT(na3168_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3168_1_i) );
// C_MX4b/D///      x99y99     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3169_1 ( .OUT(na3169_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3765_2),
                      .IN8(na9777_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3169_2 ( .OUT(na3169_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3169_1_i) );
// C_MX4b/D///      x99y108     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3170_1 ( .OUT(na3170_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9778_2),
                      .IN8(na3753_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3170_2 ( .OUT(na3170_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3170_1_i) );
// C_MX4b/D///      x115y93     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3171_1 ( .OUT(na3171_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3171_1), .IN6(na1078_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3171_2 ( .OUT(na3171_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3171_1_i) );
// C_MX4b/D///      x104y88     80'h00_FE00_00_0040_0AC3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3172_1 ( .OUT(na3172_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na261_1),
                      .IN8(na3172_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a3172_2 ( .OUT(na3172_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3172_1_i) );
// C_AND/D//AND/D      x51y114     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3173_1 ( .OUT(na3173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3809_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3173_2 ( .OUT(na3173_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3173_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3173_4 ( .OUT(na3173_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(na3809_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3173_5 ( .OUT(na3173_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3173_2_i) );
// C_MX4b/D///      x105y101     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3174_1 ( .OUT(na3174_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3174_1), .IN6(na1211_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3174_2 ( .OUT(na3174_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3174_1_i) );
// C_MX4b/D///      x120y84     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3175_1 ( .OUT(na3175_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9779_2), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3175_2 ( .OUT(na3175_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3175_1_i) );
// C_MX4b/D///      x111y58     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3177_1 ( .OUT(na3177_1_i), .IN1(~na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na6480_1), .IN6(na3177_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3177_2 ( .OUT(na3177_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3177_1_i) );
// C_///AND/D      x113y82     80'h00_FE00_80_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3178_4 ( .OUT(na3178_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na3179_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3178_5 ( .OUT(na3178_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3178_2_i) );
// C_MX2a////      x106y89     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3179_1 ( .OUT(na3179_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na9781_2), .IN4(~na159_1), .IN5(na853_2), .IN6(na459_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x115y67     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3180_1 ( .OUT(na3180_1_i), .IN1(na1728_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3180_1), .IN6(na3181_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3180_2 ( .OUT(na3180_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3180_1_i) );
// C_///AND/      x115y66     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3181_4 ( .OUT(na3181_2), .IN1(~na1730_1), .IN2(~na9782_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x49y113     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3182_1 ( .OUT(na3182_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3811_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3182_2 ( .OUT(na3182_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3182_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3182_4 ( .OUT(na3182_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3811_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3182_5 ( .OUT(na3182_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3182_2_i) );
// C_MX4b/D///      x120y99     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3183_1 ( .OUT(na3183_1_i), .IN1(na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9784_2), .IN6(na1073_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3183_2 ( .OUT(na3183_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3183_1_i) );
// C_MX4b/D///      x116y60     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3185_1 ( .OUT(na3185_1_i), .IN1(na268_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na9786_2), .IN6(na6479_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3185_2 ( .OUT(na3185_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3185_1_i) );
// C_///AND/D      x98y79     80'h00_FE00_80_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3186_4 ( .OUT(na3186_2_i), .IN1(~na3187_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3186_5 ( .OUT(na3186_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3186_2_i) );
// C_MX2a////      x97y85     80'h00_0018_00_0040_0CCC_F800
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3187_1 ( .OUT(na3187_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na3186_2), .IN4(~na159_1), .IN5(na1028_1), .IN6(na459_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x49y114     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3188_1 ( .OUT(na3188_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na971_1), .IN6(1'b1), .IN7(na3813_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3188_2 ( .OUT(na3188_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3188_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3188_4 ( .OUT(na3188_2_i), .IN1(na971_1), .IN2(1'b1), .IN3(na3813_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a3188_5 ( .OUT(na3188_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3188_2_i) );
// C_MX4b/D///      x120y100     80'h00_FE00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3189_1 ( .OUT(na3189_1_i), .IN1(~na581_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na1034_1), .IN6(na9787_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3189_2 ( .OUT(na3189_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3189_1_i) );
// C_MX4b/D///      x94y95     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3190_1 ( .OUT(na3190_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3765_1),
                      .IN8(na9788_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3190_2 ( .OUT(na3190_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3190_1_i) );
// C_MX4b/D///      x121y63     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3191_1 ( .OUT(na3191_1_i), .IN1(na444_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3191_1), .IN6(na6477_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3191_2 ( .OUT(na3191_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3191_1_i) );
// C_MX4b/D///      x100y108     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3192_1 ( .OUT(na3192_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3755_1),
                      .IN8(na3192_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3192_2 ( .OUT(na3192_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3192_1_i) );
// C_MX4b/D///      x121y89     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3193_1 ( .OUT(na3193_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3193_1), .IN6(na893_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3193_2 ( .OUT(na3193_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3193_1_i) );
// C_MX4b/D///      x107y85     80'h00_FE00_00_0040_0A3C_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3194_1 ( .OUT(na3194_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3194_1), .IN6(na262_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a3194_2 ( .OUT(na3194_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3194_1_i) );
// C_MX4b/D///      x98y97     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3195_1 ( .OUT(na3195_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3195_1),
                      .IN8(na3751_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3195_2 ( .OUT(na3195_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3195_1_i) );
// C_MX4b/D///      x121y91     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3196_1 ( .OUT(na3196_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3196_1), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3196_2 ( .OUT(na3196_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3196_1_i) );
// C_MX4b/D///      x106y92     80'h00_FE00_00_0040_0AC3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3197_1 ( .OUT(na3197_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na263_1),
                      .IN8(na3197_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a3197_2 ( .OUT(na3197_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3197_1_i) );
// C_AND/D///      x88y90     80'h00_FE00_00_0000_0888_A2AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3198_1 ( .OUT(na3198_1_i), .IN1(na4899_2), .IN2(1'b1), .IN3(na9222_2), .IN4(1'b1), .IN5(na428_2), .IN6(~na435_1), .IN7(na433_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3198_2 ( .OUT(na3198_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3198_1_i) );
// C_MX4b/D///      x86y85     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3200_1 ( .OUT(na3200_1_i), .IN1(na2680_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3200_1),
                      .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3200_2 ( .OUT(na3200_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3200_1_i) );
// C_MX4b/D///      x104y108     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3201_1 ( .OUT(na3201_1_i), .IN1(~na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3755_2),
                      .IN8(na3201_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3201_2 ( .OUT(na3201_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3201_1_i) );
// C_MX4b/D///      x117y99     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3203_1 ( .OUT(na3203_1_i), .IN1(~na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na833_1),
                      .IN8(na9790_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3203_2 ( .OUT(na3203_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3203_1_i) );
// C_AND/D///      x130y48     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3204_1 ( .OUT(na3204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3876_1), .IN6(1'b1), .IN7(1'b1), .IN8(na499_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3204_2 ( .OUT(na3204_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3204_1_i) );
// C_MX4b/D///      x103y108     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3205_1 ( .OUT(na3205_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9791_2),
                      .IN8(na3757_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3205_2 ( .OUT(na3205_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3205_1_i) );
// C_MX4b/D///      x110y92     80'h00_FE00_00_0040_0AC3_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3207_1 ( .OUT(na3207_1_i), .IN1(~na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(na264_1),
                      .IN8(na3207_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a3207_2 ( .OUT(na3207_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3207_1_i) );
// C_MX4b/D///      x95y113     80'h00_FE00_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3208_1 ( .OUT(na3208_1_i), .IN1(na248_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3208_1), .IN6(~na9792_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3208_2 ( .OUT(na3208_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3208_1_i) );
// C_MX4b/D///      x101y85     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3210_1 ( .OUT(na3210_1_i), .IN1(na448_1), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3210_1), .IN6(na265_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3210_2 ( .OUT(na3210_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3210_1_i) );
// C_MX4b/D///      x117y97     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3211_1 ( .OUT(na3211_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3211_1), .IN6(na482_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3211_2 ( .OUT(na3211_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3211_1_i) );
// C_MX4b/D///      x115y85     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3212_1 ( .OUT(na3212_1_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9793_2),
                      .IN8(na1097_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3212_2 ( .OUT(na3212_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3212_1_i) );
// C_AND////      x93y92     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3213_1 ( .OUT(na3213_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1344_2), .IN8(na1349_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x127y97     80'h00_FA18_00_0000_0888_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3214_1 ( .OUT(na3214_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2894_2), .IN7(1'b1), .IN8(na2836_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3214_5 ( .OUT(na3214_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3214_1) );
// C_OR////      x46y82     80'h00_0018_00_0000_0CEE_AE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3215_1 ( .OUT(na3215_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2867_2), .IN6(na2870_2), .IN7(na2868_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/D      x94y98     80'h00_FE00_80_0000_0C0E_FFAA
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3216_4 ( .OUT(na3216_2_i), .IN1(na3217_1), .IN2(1'b0), .IN3(na8137_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3216_5 ( .OUT(na3216_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3216_2_i) );
// C_ORAND////      x91y95     80'h00_0018_00_0000_0888_F73C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3217_1 ( .OUT(na3217_1), .IN1(1'b0), .IN2(na9795_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(~na3354_1), .IN6(~na9190_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x120y69     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3218_4 ( .OUT(na3218_2), .IN1(na900_1), .IN2(na3345_1), .IN3(na1119_1), .IN4(na1333_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D//ORAND*/D      x118y67     80'h00_FE00_80_0000_0387_3773
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3219_1 ( .OUT(na3219_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3594_1), .IN6(~na9800_2), .IN7(1'b0),
                      .IN8(~na3220_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3219_2 ( .OUT(na3219_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3219_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a3219_4 ( .OUT(na3219_2_i), .IN1(1'b0), .IN2(~na8158_1), .IN3(~na3219_2), .IN4(~na3226_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3219_5 ( .OUT(na3219_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3219_2_i) );
// C_ORAND////      x114y66     80'h00_0018_00_0000_0888_F73A
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3220_1 ( .OUT(na3220_1), .IN1(na9796_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na6626_1), .IN5(~na1730_1), .IN6(~na3343_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x119y70     80'h00_FE00_00_0000_0788_3FC7
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3222_1 ( .OUT(na3222_1_i), .IN1(~na9799_2), .IN2(~na3356_1), .IN3(1'b0), .IN4(na8142_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(~na3224_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3222_2 ( .OUT(na3222_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3222_1_i) );
// C_///AND/      x116y68     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3224_4 ( .OUT(na3224_2), .IN1(na1730_1), .IN2(na3343_1), .IN3(na3219_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y71     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3225_1 ( .OUT(na3225_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na911_2), .IN7(na1895_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x114y70     80'h00_0078_00_0000_0C88_333C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3226_1 ( .OUT(na3226_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3343_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3226_4 ( .OUT(na3226_2), .IN1(1'b1), .IN2(na3343_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x116y72     80'h00_FE00_80_0000_0C07_FF3E
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a3227_4 ( .OUT(na3227_2_i), .IN1(na3225_1), .IN2(na3228_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3227_5 ( .OUT(na3227_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3227_2_i) );
// C_ORAND////      x115y72     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3228_1 ( .OUT(na3228_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9799_2), .IN6(~na3222_1), .IN7(1'b0), .IN8(~na3227_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x45y56     80'h00_0060_00_0000_0C0E_FFEC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3229_4 ( .OUT(na3229_2), .IN1(1'b0), .IN2(na2865_2), .IN3(na2866_1), .IN4(na2863_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x59y36     80'h00_0060_00_0000_0C0E_FFEC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3230_4 ( .OUT(na3230_2), .IN1(1'b0), .IN2(na2861_1), .IN3(na2862_1), .IN4(na2863_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x45y70     80'h00_0018_00_0000_0CEE_EA00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3231_1 ( .OUT(na3231_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2860_2), .IN6(1'b0), .IN7(na2858_1), .IN8(na9702_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y97     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3232_1 ( .OUT(na3232_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1039_1), .IN6(~na6065_2), .IN7(na953_1),
                      .IN8(~na6626_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x46y64     80'h00_0060_00_0000_0C0E_FFEA
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3233_4 ( .OUT(na3233_2), .IN1(na2855_2), .IN2(1'b0), .IN3(na2857_2), .IN4(na2856_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x113y97     80'h00_0060_00_0000_0C08_FF14
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3234_4 ( .OUT(na3234_2), .IN1(~na2733_1), .IN2(na6065_2), .IN3(~na3688_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x112y92     80'h00_0018_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3237_1 ( .OUT(na3237_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8358_2), .IN6(~na6065_2), .IN7(na3238_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x120y105     80'h00_0060_00_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3238_4 ( .OUT(na3238_2), .IN1(na8154_1), .IN2(na6065_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y116     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3239_1 ( .OUT(na3239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3732_1), .IN6(na316_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y89     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3240_4 ( .OUT(na3240_2), .IN1(1'b1), .IN2(~na316_1), .IN3(na9936_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x77y90     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3241_1 ( .OUT(na3241_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2881_1), .IN7(na2882_2), .IN8(na2880_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x90y73     80'h00_0018_00_0000_0CEE_EA00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3242_1 ( .OUT(na3242_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2885_1), .IN6(1'b0), .IN7(na2882_2), .IN8(na2883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y73     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3243_1 ( .OUT(na3243_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9151_2), .IN6(1'b1), .IN7(1'b1), .IN8(na378_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x62y85     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3244_4 ( .OUT(na3244_2), .IN1(1'b1), .IN2(na2172_2), .IN3(1'b1), .IN4(na3315_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x91y48     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3247_1 ( .OUT(na3247_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2878_2), .IN7(na2876_2), .IN8(na2877_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x63y74     80'h00_0060_00_0000_0C0E_FFAE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3248_4 ( .OUT(na3248_2), .IN1(na2888_2), .IN2(na2886_2), .IN3(na2887_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x87y48     80'h00_0060_00_0000_0C0E_FFEA
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3249_4 ( .OUT(na3249_2), .IN1(na2850_2), .IN2(1'b0), .IN3(na2853_1), .IN4(na2846_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y66     80'h00_0018_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3250_1 ( .OUT(na3250_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6118_2), .IN6(na2834_1), .IN7(na2808_2),
                      .IN8(~na6626_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x109y71     80'h00_0060_00_0000_0C08_FF12
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3251_4 ( .OUT(na3251_2), .IN1(na6118_2), .IN2(~na2759_1), .IN3(~na9942_2), .IN4(~na3646_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x102y54     80'h00_0018_00_0000_0C88_DAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3253_1 ( .OUT(na3253_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6118_2), .IN6(1'b0), .IN7(~na9671_2), .IN8(na9834_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x109y60     80'h00_0060_00_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3254_4 ( .OUT(na3254_2), .IN1(na6118_2), .IN2(na8166_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y68     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3255_1 ( .OUT(na3255_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3254_2), .IN7(1'b1), .IN8(~na3253_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x117y71     80'h00_FE00_00_0000_0CEE_E000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3256_1 ( .OUT(na3256_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3257_1), .IN8(na8167_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3256_2 ( .OUT(na3256_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3256_1_i) );
// C_AND////      x116y75     80'h00_0018_00_0000_0C88_32FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3257_1 ( .OUT(na3257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3256_1), .IN6(~na3345_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////D      x117y93     80'h00_FA18_00_0000_0888_FF7C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3258_1 ( .OUT(na3258_1), .IN1(1'b0), .IN2(na2894_2), .IN3(~na2838_1), .IN4(~na2836_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3258_5 ( .OUT(na3258_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3258_1) );
// C_ORAND*/D///      x81y84     80'h00_FE00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3259_1 ( .OUT(na3259_1_i), .IN1(~na546_1), .IN2(~na9264_2), .IN3(~na531_1), .IN4(~na9751_2), .IN5(~na546_2), .IN6(~na9348_2),
                      .IN7(~na531_2), .IN8(~na1175_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3259_2 ( .OUT(na3259_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3259_1_i) );
// C_AND/D///      x69y75     80'h00_FA00_00_0000_0C88_83FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3262_1 ( .OUT(na3262_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na365_2), .IN7(na2558_1), .IN8(na2556_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3262_2 ( .OUT(na3262_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3262_1_i) );
// C_MX2a/D///      x55y62     80'h00_FA00_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3263_1 ( .OUT(na3263_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na2558_1), .IN4(na8173_1), .IN5(~na2555_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3263_2 ( .OUT(na3263_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3263_1_i) );
// C_MX2a/D///      x57y73     80'h00_FA00_00_0040_0C0A_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3264_1 ( .OUT(na3264_1_i), .IN1(1'b0), .IN2(na2554_1), .IN3(1'b0), .IN4(na8174_2), .IN5(1'b1), .IN6(1'b1), .IN7(na2558_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3264_2 ( .OUT(na3264_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3264_1_i) );
// C_MX2a/D///      x62y75     80'h00_FA00_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3265_1 ( .OUT(na3265_1_i), .IN1(1'b0), .IN2(na2554_1), .IN3(1'b0), .IN4(na8175_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2556_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3265_2 ( .OUT(na3265_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3265_1_i) );
// C_ORAND/D///      x46y85     80'h00_FA00_00_0000_0888_FAE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3266_1 ( .OUT(na3266_1_i), .IN1(1'b0), .IN2(~na2554_1), .IN3(na8176_1), .IN4(na9623_2), .IN5(na2566_1), .IN6(1'b0), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3266_2 ( .OUT(na3266_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3266_1_i) );
// C_///OR/D      x52y45     80'h00_FA00_80_0000_0C0E_FFAC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3268_4 ( .OUT(na3268_2_i), .IN1(1'b0), .IN2(na2554_1), .IN3(na8177_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3268_5 ( .OUT(na3268_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3268_2_i) );
// C_///ORAND*/D      x69y77     80'h00_FA00_80_0000_0C07_FFDB
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a3269_4 ( .OUT(na3269_2_i), .IN1(na2566_1), .IN2(~na2564_1), .IN3(~na9622_2), .IN4(na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3269_5 ( .OUT(na3269_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3269_2_i) );
// C_ORAND/D///      x75y78     80'h00_FA00_00_0000_0888_C35D
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3270_1 ( .OUT(na3270_1_i), .IN1(~na2566_1), .IN2(na9626_2), .IN3(~na2558_1), .IN4(1'b0), .IN5(1'b0), .IN6(~na2554_1), .IN7(1'b0),
                      .IN8(na3272_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3270_2 ( .OUT(na3270_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3270_1_i) );
// C_///AND/      x70y80     80'h00_0060_00_0000_0C08_FFC4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3272_4 ( .OUT(na3272_2), .IN1(~na2565_1), .IN2(na2564_1), .IN3(1'b1), .IN4(na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x72y94     80'h00_0018_00_0000_0CEE_EA00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3273_1 ( .OUT(na3273_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2839_1), .IN6(1'b0), .IN7(na2844_2), .IN8(na2846_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y76     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3274_4 ( .OUT(na3274_2), .IN1(na6118_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1425_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y41     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3275_1 ( .OUT(na3275_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3664_1), .IN8(na1425_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x98y101     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3276_1 ( .OUT(na3276_1_i), .IN1(na3354_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(na3276_1),
                      .IN8(na9814_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3276_2 ( .OUT(na3276_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3276_1_i) );
// C_AND////      x91y98     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3277_1 ( .OUT(na3277_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na279_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na272_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x96y99     80'h00_0060_00_0000_0C0E_FF5C
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3278_4 ( .OUT(na3278_2), .IN1(1'b0), .IN2(na8182_1), .IN3(~na3279_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x88y85     80'h00_0018_00_0040_0CF9_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3279_1 ( .OUT(na3279_1), .IN1(~na5451_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na5450_1), .IN5(~na279_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na272_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x49y84     80'h00_0018_00_0040_0C99_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3280_1 ( .OUT(na3280_1), .IN1(~na2389_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na3281_1), .IN5(~na3326_2), .IN6(1'b1), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y72     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3281_1 ( .OUT(na3281_1), .IN1(~na50_1), .IN2(1'b1), .IN3(~na357_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x114y69     80'h00_0018_00_0000_0CEE_A300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3282_1 ( .OUT(na3282_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3283_1), .IN7(na8185_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x113y68     80'h00_0018_00_0040_0CF6_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3283_1 ( .OUT(na3283_1), .IN1(1'b1), .IN2(~na5216_2), .IN3(~na5217_1), .IN4(1'b1), .IN5(na3180_1), .IN6(1'b1), .IN7(na2163_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y66     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3284_4 ( .OUT(na3284_2), .IN1(~na3180_1), .IN2(1'b1), .IN3(~na2163_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x109y65     80'h00_0018_00_0000_0CEE_C300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3285_1 ( .OUT(na3285_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3286_1), .IN7(1'b0), .IN8(na8186_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x113y72     80'h00_0018_00_0040_0CF6_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3286_1 ( .OUT(na3286_1), .IN1(1'b1), .IN2(~na5220_1), .IN3(~na5221_2), .IN4(1'b1), .IN5(na3180_1), .IN6(1'b1), .IN7(na2163_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x95y99     80'h00_0060_00_0000_0C0E_FF3C
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3287_4 ( .OUT(na3287_2), .IN1(1'b0), .IN2(na8187_1), .IN3(1'b0), .IN4(~na3288_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x94y92     80'h00_0018_00_0040_0CF6_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3288_1 ( .OUT(na3288_1), .IN1(1'b1), .IN2(~na5447_1), .IN3(~na5446_2), .IN4(1'b1), .IN5(na279_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na272_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x87y66     80'h00_0060_00_0000_0C0E_FFAE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3289_4 ( .OUT(na3289_2), .IN1(na2872_1), .IN2(na2870_2), .IN3(na2871_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x113y73     80'h00_FE00_00_0000_0788_3FB7
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3290_1 ( .OUT(na3290_1_i), .IN1(~na9831_2), .IN2(~na3345_1), .IN3(na4204_2), .IN4(~na9811_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(~na6626_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3290_2 ( .OUT(na3290_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3290_1_i) );
// C_ORAND*/D///      x94y119     80'h00_FE00_00_0000_0788_7F33
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3292_1 ( .OUT(na3292_1_i), .IN1(1'b0), .IN2(~na8190_2), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3357_1),
                      .IN8(~na9832_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3292_2 ( .OUT(na3292_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3292_1_i) );
// C_ORAND////      x93y120     80'h00_0018_00_0000_0888_7F3A
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3296_1 ( .OUT(na3296_1), .IN1(na3297_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3357_1),
                      .IN8(~na9195_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D//OR/D      x91y119     80'h00_FE00_80_0000_0CEE_CA0E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3297_1 ( .OUT(na3297_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na8192_2), .IN6(1'b0), .IN7(1'b0), .IN8(na3298_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3297_2 ( .OUT(na3297_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3297_1_i) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3297_4 ( .OUT(na3297_2_i), .IN1(na8192_1), .IN2(na3296_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3297_5 ( .OUT(na3297_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3297_2_i) );
// C_AND////      x100y98     80'h00_0018_00_0000_0C88_1AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3298_1 ( .OUT(na3298_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3297_1), .IN6(1'b1), .IN7(~na3357_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x97y94     80'h00_FE00_80_0000_0C07_FF3E
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a3299_4 ( .OUT(na3299_2_i), .IN1(na3300_2), .IN2(na3213_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3299_5 ( .OUT(na3299_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3299_2_i) );
// C_///ORAND/      x89y91     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3300_4 ( .OUT(na3300_2), .IN1(~na3354_1), .IN2(~na9828_2), .IN3(~na9813_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y99     80'h00_FE00_00_0000_0CEE_CC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3301_1 ( .OUT(na3301_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3302_1), .IN7(1'b0), .IN8(na8197_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3301_2 ( .OUT(na3301_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3301_1_i) );
// C_ORAND////      x85y90     80'h00_0018_00_0000_0888_FE3C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3302_1 ( .OUT(na3302_1), .IN1(1'b0), .IN2(na3213_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(na3588_1), .IN6(na3299_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x63y38     80'h00_0018_00_0000_0CEE_CE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3303_1 ( .OUT(na3303_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2888_2), .IN6(na2891_2), .IN7(1'b0), .IN8(na2890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x91y52     80'h00_0060_00_0000_0C0E_FFAE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3304_4 ( .OUT(na3304_2), .IN1(na2875_1), .IN2(na2873_1), .IN3(na2876_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x79y83     80'h00_FA00_00_0000_0888_8284
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3305_1 ( .OUT(na3305_1_i), .IN1(~na2584_2), .IN2(na9624_2), .IN3(na3307_1), .IN4(na2572_1), .IN5(na2569_1), .IN6(~na2586_2),
                      .IN7(na3307_2), .IN8(na389_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3305_2 ( .OUT(na3305_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3305_1_i) );
// C_AND///AND/      x80y93     80'h00_0078_00_0000_0C88_C833
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3307_1 ( .OUT(na3307_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2570_1), .IN6(na2571_1), .IN7(1'b1), .IN8(na2573_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3307_4 ( .OUT(na3307_2), .IN1(1'b1), .IN2(~na2567_1), .IN3(1'b1), .IN4(~na2592_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x70y111     80'h00_FA00_00_0000_0888_8224
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3308_1 ( .OUT(na3308_1_i), .IN1(~na2584_2), .IN2(na9624_2), .IN3(na3307_1), .IN4(~na2572_1), .IN5(na2569_1), .IN6(~na2586_2),
                      .IN7(na3307_2), .IN8(na389_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3308_2 ( .OUT(na3308_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3308_1_i) );
// C_AND/D//AND/D      x66y110     80'h00_FA00_80_0000_0C88_8881
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3309_1 ( .OUT(na3309_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2584_2), .IN6(na2586_2), .IN7(na3311_1),
                      .IN8(na389_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3309_2 ( .OUT(na3309_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3309_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3309_4 ( .OUT(na3309_2_i), .IN1(~na2584_2), .IN2(~na2586_2), .IN3(na3316_1), .IN4(na389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3309_5 ( .OUT(na3309_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3309_2_i) );
// C_AND////      x78y95     80'h00_0018_00_0000_0888_242A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3311_1 ( .OUT(na3311_1), .IN1(na2570_1), .IN2(1'b1), .IN3(na3307_2), .IN4(~na2573_1), .IN5(~na2569_1), .IN6(na2571_1), .IN7(na2568_1),
                      .IN8(~na2572_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x59y111     80'h00_FA00_80_0000_0C88_8482
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3313_1 ( .OUT(na3313_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2584_2), .IN6(na2586_2), .IN7(na3311_1),
                      .IN8(na389_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3313_2 ( .OUT(na3313_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3313_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3313_4 ( .OUT(na3313_2_i), .IN1(na2584_2), .IN2(~na2586_2), .IN3(na3311_1), .IN4(na389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3313_5 ( .OUT(na3313_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3313_2_i) );
// C_AND/D///      x80y94     80'h00_FA00_00_0000_0888_AF22
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3315_1 ( .OUT(na3315_1_i), .IN1(na2584_2), .IN2(~na2586_2), .IN3(na2588_2), .IN4(~na2590_2), .IN5(1'b1), .IN6(1'b1), .IN7(na3316_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3315_2 ( .OUT(na3315_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3315_1_i) );
// C_AND////      x80y89     80'h00_0018_00_0000_0888_142A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3316_1 ( .OUT(na3316_1), .IN1(na2570_1), .IN2(1'b1), .IN3(na3307_2), .IN4(~na2573_1), .IN5(~na2569_1), .IN6(na2571_1), .IN7(~na2568_1),
                      .IN8(~na2572_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x71y100     80'h00_FA00_00_0000_0888_A523
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3317_1 ( .OUT(na3317_1_i), .IN1(1'b1), .IN2(~na2586_2), .IN3(na2588_2), .IN4(~na2590_2), .IN5(~na2584_2), .IN6(1'b1), .IN7(na3316_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3317_2 ( .OUT(na3317_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3317_1_i) );
// C_AND/D///      x80y100     80'h00_FA00_00_0000_0888_A523
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3319_1 ( .OUT(na3319_1_i), .IN1(1'b1), .IN2(~na2586_2), .IN3(na2588_2), .IN4(~na2590_2), .IN5(~na2584_2), .IN6(1'b1), .IN7(na3311_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3319_2 ( .OUT(na3319_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3319_1_i) );
// C_AND/D///      x80y85     80'h00_FA00_00_0000_0C88_84FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3321_1 ( .OUT(na3321_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2570_1), .IN6(na365_2), .IN7(na2558_1),
                      .IN8(na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3321_2 ( .OUT(na3321_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3321_1_i) );
// C_AND/D///      x80y84     80'h00_FA00_00_0000_0888_4FA8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3323_1 ( .OUT(na3323_1_i), .IN1(na2570_1), .IN2(na365_2), .IN3(na2558_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2588_2),
                      .IN8(na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3323_2 ( .OUT(na3323_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3323_1_i) );
// C_AND*/D///      x72y82     80'h00_FA00_00_0000_0788_2531
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a3324_1 ( .OUT(na3324_1_i), .IN1(~na2576_2), .IN2(~na2578_2), .IN3(1'b1), .IN4(~na2580_2), .IN5(~na2574_2), .IN6(1'b1), .IN7(na9622_2),
                      .IN8(~na2582_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3324_2 ( .OUT(na3324_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3324_1_i) );
// C_AND/D///      x77y74     80'h00_FA00_00_0000_0C88_15FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3325_1 ( .OUT(na3325_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2555_1), .IN6(1'b1), .IN7(~na2558_1),
                      .IN8(~na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3325_2 ( .OUT(na3325_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3325_1_i) );
// C_///AND/D      x55y77     80'h00_FA00_80_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3326_4 ( .OUT(na3326_2_i), .IN1(~na2566_1), .IN2(~na2554_1), .IN3(na9622_2), .IN4(na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3326_5 ( .OUT(na3326_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3326_2_i) );
// C_///AND/D      x83y77     80'h00_FA00_80_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3327_4 ( .OUT(na3327_2_i), .IN1(na2565_1), .IN2(~na2564_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3327_5 ( .OUT(na3327_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3327_2_i) );
// C_AND/D///      x69y73     80'h00_FA00_00_0000_0C88_42FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3328_1 ( .OUT(na3328_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2566_1), .IN6(~na2554_1), .IN7(~na2558_1),
                      .IN8(na3272_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3328_2 ( .OUT(na3328_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3328_1_i) );
// C_///AND/D      x59y61     80'h00_FA00_80_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3329_4 ( .OUT(na3329_2_i), .IN1(~na2555_1), .IN2(1'b1), .IN3(na2558_1), .IN4(~na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3329_5 ( .OUT(na3329_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3329_2_i) );
// C_ORAND/D///      x63y74     80'h00_FA00_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3330_1 ( .OUT(na3330_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8362_2), .IN6(na2554_1), .IN7(~na3331_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3330_2 ( .OUT(na3330_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3330_1_i) );
// C_MX4b////      x76y67     80'h00_0018_00_0040_0A3F_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3331_1 ( .OUT(na3331_1), .IN1(1'b1), .IN2(na2554_1), .IN3(na2558_1), .IN4(1'b1), .IN5(~na9808_2), .IN6(~na2557_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x63y70     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3332_1 ( .OUT(na3332_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3328_1), .IN6(na3270_1), .IN7(1'b1), .IN8(na2421_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////D      x118y103     80'h00_FE18_00_0000_0888_FF6A
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3333_1 ( .OUT(na3333_1), .IN1(~na951_1), .IN2(1'b0), .IN3(na9387_2), .IN4(~na9389_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3333_5 ( .OUT(na3333_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3333_1) );
// C_///AND/      x46y93     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3334_4 ( .OUT(na3334_2), .IN1(na9943_2), .IN2(na6665_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x75y97     80'h00_0060_00_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3335_4 ( .OUT(na3335_2), .IN1(na402_1), .IN2(na401_2), .IN3(1'b0), .IN4(~na341_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x75y93     80'h00_0018_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3337_1 ( .OUT(na3337_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na402_1), .IN6(na401_2), .IN7(1'b0), .IN8(~na378_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x117y78     80'h00_0060_00_0000_0C08_FFA4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3339_4 ( .OUT(na3339_2), .IN1(~na1020_1), .IN2(na1012_1), .IN3(na1021_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x113y100     80'h00_0018_00_0000_0C88_A4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3340_1 ( .OUT(na3340_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1006_2), .IN6(na1007_1), .IN7(na997_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x117y96     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3341_1 ( .OUT(na3341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1006_2), .IN6(na1007_1), .IN7(na997_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y68     80'h00_0018_00_0000_0888_58F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3342_1 ( .OUT(na3342_1), .IN1(~na3594_1), .IN2(~na3356_1), .IN3(1'b1), .IN4(1'b1), .IN5(na3225_1), .IN6(na3555_1), .IN7(~na3219_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x121y62     80'h00_FE00_00_0000_0888_F1C2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3343_1 ( .OUT(na3343_1_i), .IN1(na985_2), .IN2(~na2972_1), .IN3(1'b1), .IN4(na500_2), .IN5(~na985_1), .IN6(~na2972_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3343_2 ( .OUT(na3343_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3343_1_i) );
// C_AND/D///      x121y70     80'h00_FE00_00_0000_0888_F483
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3345_1 ( .OUT(na3345_1_i), .IN1(1'b1), .IN2(~na2718_1), .IN3(na2737_1), .IN4(na500_2), .IN5(~na2746_2), .IN6(na2718_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3345_2 ( .OUT(na3345_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3345_1_i) );
// C_///AND/      x107y92     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3347_4 ( .OUT(na3347_2), .IN1(~na1006_2), .IN2(~na1007_1), .IN3(na997_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y76     80'h00_0018_00_0000_0C88_54FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3348_1 ( .OUT(na3348_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1020_1), .IN6(na1012_1), .IN7(~na1021_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y76     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3349_4 ( .OUT(na3349_2), .IN1(na1020_1), .IN2(na1012_1), .IN3(na1021_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x114y76     80'h00_0018_00_0000_0C88_58FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3350_1 ( .OUT(na3350_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1020_1), .IN6(na1012_1), .IN7(~na1021_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x107y96     80'h00_0060_00_0000_0C08_FFA2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3351_4 ( .OUT(na3351_2), .IN1(na1006_2), .IN2(~na1007_1), .IN3(na997_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x111y73     80'h00_FE00_80_0000_0C08_FF32
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3352_4 ( .OUT(na3352_2_i), .IN1(na3352_2), .IN2(~na3345_1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3352_5 ( .OUT(na3352_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3352_2_i) );
// C_ORAND////      x98y92     80'h00_0018_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3353_1 ( .OUT(na3353_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na285_1), .IN6(~na7348_1), .IN7(na9794_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x91y103     80'h00_FE00_00_0000_0888_5C43
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3354_1 ( .OUT(na3354_1_i), .IN1(1'b1), .IN2(~na291_1), .IN3(~na289_1), .IN4(na325_2), .IN5(1'b1), .IN6(na291_2), .IN7(~na289_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3354_2 ( .OUT(na3354_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3354_1_i) );
// C_AND/D///      x115y68     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3356_1 ( .OUT(na3356_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3356_1), .IN7(1'b1), .IN8(na3226_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3356_2 ( .OUT(na3356_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3356_1_i) );
// C_AND/D///      x96y103     80'h00_FE00_00_0000_0888_A54C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3357_1 ( .OUT(na3357_1_i), .IN1(1'b1), .IN2(na334_1), .IN3(~na336_1), .IN4(na325_2), .IN5(~na338_2), .IN6(1'b1), .IN7(na336_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3357_2 ( .OUT(na3357_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3357_1_i) );
// C_///AND/      x58y78     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3359_4 ( .OUT(na3359_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(na3266_1), .IN4(~na3360_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y74     80'h00_0018_00_0040_0AB4_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3360_1 ( .OUT(na3360_1), .IN1(~na50_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na355_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y84     80'h00_0018_00_0000_0C88_45FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3361_1 ( .OUT(na3361_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(~na3362_1), .IN8(na9805_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y73     80'h00_0018_00_0040_0AB4_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3362_1 ( .OUT(na3362_1), .IN1(1'b1), .IN2(~na9826_2), .IN3(1'b1), .IN4(~na9254_2), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y84     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3363_1 ( .OUT(na3363_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(na3266_1), .IN8(~na3364_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y76     80'h00_0018_00_0040_0AB4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3364_1 ( .OUT(na3364_1), .IN1(1'b1), .IN2(~na3489_1), .IN3(~na545_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y81     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3365_4 ( .OUT(na3365_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(na3266_1), .IN4(~na3366_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y74     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3366_1 ( .OUT(na3366_1), .IN1(~na3487_1), .IN2(1'b1), .IN3(~na550_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y81     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3367_1 ( .OUT(na3367_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3368_1), .IN6(~na9819_2), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y69     80'h00_0018_00_0040_0AB4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3368_1 ( .OUT(na3368_1), .IN1(1'b1), .IN2(~na9593_2), .IN3(~na2369_2), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x47y82     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3369_4 ( .OUT(na3369_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(na3266_1), .IN4(~na3370_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y68     80'h00_0018_00_0040_0AB4_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3370_1 ( .OUT(na3370_1), .IN1(~na2362_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2348_2), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x46y84     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3371_4 ( .OUT(na3371_2), .IN1(~na3326_2), .IN2(~na3372_1), .IN3(na3266_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y78     80'h00_0018_00_0040_0AB4_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3372_1 ( .OUT(na3372_1), .IN1(na2309_2), .IN2(1'b1), .IN3(na589_2), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y83     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3373_1 ( .OUT(na3373_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(na3266_1), .IN8(~na3374_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y72     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3374_1 ( .OUT(na3374_1), .IN1(~na2338_2), .IN2(1'b1), .IN3(~na589_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y84     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3375_4 ( .OUT(na3375_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(na3266_1), .IN4(~na3376_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y76     80'h00_0018_00_0040_0AB4_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3376_1 ( .OUT(na3376_1), .IN1(1'b1), .IN2(~na9581_2), .IN3(1'b1), .IN4(~na594_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y84     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3377_1 ( .OUT(na3377_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(~na3378_1), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y72     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3378_1 ( .OUT(na3378_1), .IN1(~na2332_2), .IN2(1'b1), .IN3(~na2327_2), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x47y84     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3379_4 ( .OUT(na3379_2), .IN1(~na3326_2), .IN2(~na3380_1), .IN3(na3266_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y72     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3380_1 ( .OUT(na3380_1), .IN1(~na2378_2), .IN2(1'b1), .IN3(~na2316_2), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x47y83     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3381_4 ( .OUT(na3381_2), .IN1(~na3326_2), .IN2(~na3382_1), .IN3(na3266_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y76     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3382_1 ( .OUT(na3382_1), .IN1(~na2378_1), .IN2(1'b1), .IN3(~na607_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y85     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3383_1 ( .OUT(na3383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(~na3384_1), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y74     80'h00_0018_00_0040_0AB4_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3384_1 ( .OUT(na3384_1), .IN1(~na9586_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na612_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x43y86     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3385_4 ( .OUT(na3385_2), .IN1(~na3326_2), .IN2(~na3386_1), .IN3(na3266_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y78     80'h00_0018_00_0040_0AB4_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3386_1 ( .OUT(na3386_1), .IN1(~na2354_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na622_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x47y82     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3387_1 ( .OUT(na3387_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(na3266_1), .IN8(~na3388_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y70     80'h00_0018_00_0040_0AB4_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3388_1 ( .OUT(na3388_1), .IN1(~na2383_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na617_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x47y83     80'h00_0018_00_0000_0C88_45FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3389_1 ( .OUT(na3389_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(~na3390_1), .IN8(na9805_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y71     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3390_1 ( .OUT(na3390_1), .IN1(~na2383_1), .IN2(1'b1), .IN3(~na627_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x47y85     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3391_4 ( .OUT(na3391_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(na3266_1), .IN4(~na3392_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y78     80'h00_0018_00_0040_0AB4_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3392_1 ( .OUT(na3392_1), .IN1(na1603_1), .IN2(1'b1), .IN3(na2369_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y85     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3393_1 ( .OUT(na3393_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(~na3394_1), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y74     80'h00_0018_00_0040_0AB4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3394_1 ( .OUT(na3394_1), .IN1(1'b1), .IN2(~na9591_2), .IN3(~na632_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y86     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3395_1 ( .OUT(na3395_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(na3266_1), .IN8(~na3396_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y76     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3396_1 ( .OUT(na3396_1), .IN1(~na2332_1), .IN2(1'b1), .IN3(~na637_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y86     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3397_1 ( .OUT(na3397_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(na3266_1), .IN8(~na3398_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y74     80'h00_0018_00_0040_0AB4_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3398_1 ( .OUT(na3398_1), .IN1(na1586_1), .IN2(1'b1), .IN3(na2357_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y89     80'h00_0018_00_0000_0C88_45FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3399_1 ( .OUT(na3399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(~na3400_1), .IN8(na9805_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y75     80'h00_0018_00_0040_0AB4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3400_1 ( .OUT(na3400_1), .IN1(1'b1), .IN2(~na2314_2), .IN3(~na661_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y91     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3401_1 ( .OUT(na3401_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(~na3402_1), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y80     80'h00_0018_00_0040_0AB4_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3402_1 ( .OUT(na3402_1), .IN1(1'b1), .IN2(~na9572_2), .IN3(1'b1), .IN4(~na667_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y84     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3403_4 ( .OUT(na3403_2), .IN1(~na3326_2), .IN2(~na3404_1), .IN3(na3266_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y80     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3404_1 ( .OUT(na3404_1), .IN1(~na2351_2), .IN2(1'b1), .IN3(~na672_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y88     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3405_1 ( .OUT(na3405_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(~na3406_1), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y80     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3406_1 ( .OUT(na3406_1), .IN1(~na9584_2), .IN2(1'b1), .IN3(~na677_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y87     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3407_4 ( .OUT(na3407_2), .IN1(~na3326_2), .IN2(~na3408_1), .IN3(na3266_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y78     80'h00_0018_00_0040_0AB4_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3408_1 ( .OUT(na3408_1), .IN1(1'b1), .IN2(~na2340_2), .IN3(1'b1), .IN4(~na682_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y85     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3409_4 ( .OUT(na3409_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(na3266_1), .IN4(~na3410_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y80     80'h00_0018_00_0040_0AB4_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3410_1 ( .OUT(na3410_1), .IN1(1'b1), .IN2(~na9576_2), .IN3(1'b1), .IN4(~na9311_2), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y88     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3411_1 ( .OUT(na3411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(~na3412_1), .IN7(na3266_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y80     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3412_1 ( .OUT(na3412_1), .IN1(~na9569_2), .IN2(1'b1), .IN3(~na692_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y88     80'h00_0060_00_0000_0C08_FF45
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3413_4 ( .OUT(na3413_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(~na3414_1), .IN4(na9805_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y79     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3414_1 ( .OUT(na3414_1), .IN1(~na2309_1), .IN2(1'b1), .IN3(~na9315_2), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y87     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3415_1 ( .OUT(na3415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3326_2), .IN6(1'b1), .IN7(na3266_1), .IN8(~na3416_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y80     80'h00_0018_00_0040_0AB4_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3416_1 ( .OUT(na3416_1), .IN1(~na2385_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na702_1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x47y86     80'h00_0060_00_0000_0C08_FF45
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3417_4 ( .OUT(na3417_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(~na3418_1), .IN4(na9805_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y77     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3418_1 ( .OUT(na3418_1), .IN1(~na2351_1), .IN2(1'b1), .IN3(~na707_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y88     80'h00_0060_00_0000_0C08_FF25
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3419_4 ( .OUT(na3419_2), .IN1(~na3326_2), .IN2(1'b1), .IN3(na3266_1), .IN4(~na3420_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y78     80'h00_0018_00_0040_0AB4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3420_1 ( .OUT(na3420_1), .IN1(~na2354_2), .IN2(1'b1), .IN3(~na723_1), .IN4(1'b1), .IN5(na10035_2), .IN6(na8184_2), .IN7(1'b1),
                      .IN8(na8183_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x75y107     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3421_1 ( .OUT(na3421_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3335_2), .IN6(~na713_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x96y100     80'h00_FE00_00_0000_0C88_45FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3423_1 ( .OUT(na3423_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9940_2), .IN6(1'b1), .IN7(~na3357_1),
                      .IN8(na3423_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3423_2 ( .OUT(na3423_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3423_1_i) );
// C_///AND/D      x91y98     80'h00_FE00_80_0000_0C08_FF34
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3424_4 ( .OUT(na3424_2_i), .IN1(~na3354_1), .IN2(na3424_2), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3424_5 ( .OUT(na3424_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3424_2_i) );
// C_MX4a////      x53y56     80'h00_0018_00_0040_0CEC_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3486_1 ( .OUT(na3486_1), .IN1(1'b0), .IN2(1'b1), .IN3(~na5965_2), .IN4(~na6310_1), .IN5(1'b1), .IN6(na369_2), .IN7(na3268_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y63     80'h00_0018_00_0040_0ACD_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3487_1 ( .OUT(na3487_1), .IN1(1'b1), .IN2(~na3486_1), .IN3(~na3268_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b0), .IN7(~na5965_1),
                      .IN8(~na5232_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x53y63     80'h00_0018_00_0040_0CEC_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3488_1 ( .OUT(na3488_1), .IN1(1'b0), .IN2(1'b1), .IN3(~na5964_2), .IN4(~na6309_2), .IN5(1'b1), .IN6(na369_2), .IN7(na3268_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y68     80'h00_0018_00_0040_0ACD_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3489_1 ( .OUT(na3489_1), .IN1(~na3488_1), .IN2(1'b1), .IN3(~na3268_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b0), .IN7(~na5964_1),
                      .IN8(~na5231_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x51y57     80'h00_0018_00_0040_0CB3_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3490_1 ( .OUT(na3490_1), .IN1(~na5963_2), .IN2(~na9937_2), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(na369_2), .IN7(~na3268_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y61     80'h00_0018_00_0040_0A37_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3491_1 ( .OUT(na3491_1), .IN1(~na3490_1), .IN2(1'b1), .IN3(na3268_2), .IN4(1'b1), .IN5(~na5963_1), .IN6(~na9866_2), .IN7(1'b1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x100y82     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3492_1 ( .OUT(na3492_1), .IN1(1'b1), .IN2(na99_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na100_2), .IN6(~na8267_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x121y107     80'h00_FA18_00_0000_0788_7F7D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3494_1 ( .OUT(na3494_1), .IN1(~na103_1), .IN2(na8271_1), .IN3(~na102_1), .IN4(~na3492_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na106_1),
                      .IN8(~na6467_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3494_5 ( .OUT(na3494_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3494_1) );
// C_ORAND*////D      x123y103     80'h00_FA18_00_0000_0788_DF7D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3496_1 ( .OUT(na3496_1), .IN1(~na103_1), .IN2(na8274_2), .IN3(~na106_1), .IN4(~na6470_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na106_2),
                      .IN8(na125_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3496_5 ( .OUT(na3496_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3496_1) );
// C_MX4a////      x91y85     80'h00_0018_00_0040_0CBA_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3497_1 ( .OUT(na3497_1), .IN1(1'b1), .IN2(~na2965_1), .IN3(1'b0), .IN4(~na796_1), .IN5(1'b1), .IN6(na2935_1), .IN7(~na2937_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x96y94     80'h00_0018_00_0040_0A3B_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3498_1 ( .OUT(na3498_1), .IN1(na3497_1), .IN2(1'b1), .IN3(1'b1), .IN4(na9714_2), .IN5(~na2963_1), .IN6(~na2964_1), .IN7(1'b0),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x114y98     80'h00_FA18_00_0000_0888_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3499_1 ( .OUT(na3499_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na103_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3498_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3499_5 ( .OUT(na3499_2), .CLK(na4116_1), .EN(na3347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3499_1) );
// C_OR////      x53y41     80'h00_0018_00_0000_0EEE_D537
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3501_1 ( .OUT(na3501_1), .IN1(~na8275_2), .IN2(~na6812_1), .IN3(1'b0), .IN4(~na8277_2), .IN5(~na8275_1), .IN6(1'b0), .IN7(~na1387_1),
                      .IN8(na8277_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x56y36     80'h00_0018_00_0000_0EEE_3C77
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3503_1 ( .OUT(na3503_1), .IN1(~na6805_1), .IN2(~na8280_2), .IN3(~na1387_1), .IN4(~na8278_2), .IN5(1'b0), .IN6(na8280_1),
                      .IN7(1'b0), .IN8(~na8278_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x74y81     80'h00_0018_00_0000_0CEE_BE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3504_1 ( .OUT(na3504_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3508_1), .IN6(na3512_1), .IN7(na3514_1),
                      .IN8(~na3503_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y53     80'h00_0018_00_0000_0888_8A88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3508_1 ( .OUT(na3508_1), .IN1(na10049_2), .IN2(na1383_1), .IN3(na8285_1), .IN4(na8283_1), .IN5(na8286_2), .IN6(1'b1), .IN7(na517_1),
                      .IN8(na8283_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x53y40     80'h00_0018_00_0000_0888_8C88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3512_1 ( .OUT(na3512_1), .IN1(na1372_1), .IN2(na8289_1), .IN3(na1387_2), .IN4(na8288_1), .IN5(1'b1), .IN6(na8289_2), .IN7(na8287_1),
                      .IN8(na10050_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x58y45     80'h00_0018_00_0000_0888_88C8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3514_1 ( .OUT(na3514_1), .IN1(na6807_2), .IN2(na5985_1), .IN3(1'b1), .IN4(na8294_1), .IN5(na10051_2), .IN6(na8292_1), .IN7(na517_2),
                      .IN8(na8294_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y55     80'h00_0018_00_0000_0888_888C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3521_1 ( .OUT(na3521_1), .IN1(1'b1), .IN2(na5985_1), .IN3(na8304_1), .IN4(na9248_2), .IN5(na8305_1), .IN6(na10052_2), .IN7(na8304_2),
                      .IN8(na8302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y68     80'h00_0018_00_0000_0888_88C8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3525_1 ( .OUT(na3525_1), .IN1(na8307_1), .IN2(na1383_1), .IN3(1'b1), .IN4(na8309_2), .IN5(na8307_2), .IN6(na8310_2), .IN7(na517_1),
                      .IN8(na8309_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x76y66     80'h00_0018_00_0000_0EEE_7BBE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3526_1 ( .OUT(na3526_1), .IN1(na2559_1), .IN2(na9629_2), .IN3(na2568_1), .IN4(~na3607_1), .IN5(na2569_1), .IN6(~na383_2),
                      .IN7(~na386_1), .IN8(~na385_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y82     80'h00_0018_00_0040_0AFD_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3527_1 ( .OUT(na3527_1), .IN1(na2566_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2556_1), .IN5(~na2565_1), .IN6(na9618_2), .IN7(~na2558_1),
                      .IN8(~na9619_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x77y78     80'h00_0018_00_0000_0888_5111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3529_1 ( .OUT(na3529_1), .IN1(~na2569_1), .IN2(~na2571_1), .IN3(~na8312_1), .IN4(~na2573_1), .IN5(~na2570_1), .IN6(~na2567_1),
                      .IN7(~na2568_1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x82y69     80'h00_0018_00_0040_0C29_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3530_1 ( .OUT(na3530_1), .IN1(na2565_1), .IN2(1'b1), .IN3(1'b0), .IN4(na8313_2), .IN5(1'b1), .IN6(na2564_1), .IN7(~na2558_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x77y71     80'h00_0018_00_0040_0CA5_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3531_1 ( .OUT(na3531_1), .IN1(na8314_1), .IN2(1'b1), .IN3(na2558_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2554_1), .IN7(~na3530_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x74y66     80'h00_0018_00_0040_0C0B_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3532_1 ( .OUT(na3532_1), .IN1(na9616_2), .IN2(na8315_2), .IN3(1'b0), .IN4(na2556_1), .IN5(na3531_1), .IN6(1'b1), .IN7(~na2558_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y65     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3535_1 ( .OUT(na3535_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na2558_1), .IN4(1'b1), .IN5(1'b0), .IN6(na2557_1), .IN7(1'b0), .IN8(na8318_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x71y87     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3537_1 ( .OUT(na3537_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na546_1), .IN6(1'b0), .IN7(na3308_1), .IN8(na8322_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x70y114     80'h00_0018_00_0000_0888_8431
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3539_1 ( .OUT(na3539_1), .IN1(~na6870_1), .IN2(~na8324_2), .IN3(1'b1), .IN4(~na6868_2), .IN5(~na3537_1), .IN6(na6869_2),
                      .IN7(na6867_1), .IN8(na8323_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x136y80     80'h00_0018_00_0040_0A8E_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3540_1 ( .OUT(na3540_1), .IN1(1'b1), .IN2(~na2894_2), .IN3(1'b1), .IN4(~na2836_2), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(~na8325_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x129y77     80'h00_0018_00_0000_0888_131F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3542_1 ( .OUT(na3542_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na298_2), .IN4(~na649_2), .IN5(1'b1), .IN6(~na8327_1), .IN7(~na298_1),
                      .IN8(~na92_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x136y84     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3543_1 ( .OUT(na3543_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2838_1), .IN8(na2836_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x126y73     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3544_1 ( .OUT(na3544_1), .IN1(1'b1), .IN2(na9697_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8328_2), .IN8(~na655_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y75     80'h00_0018_00_0000_0888_154F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3546_1 ( .OUT(na3546_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na298_1), .IN4(na8329_1), .IN5(~na214_1), .IN6(1'b1), .IN7(~na656_1),
                      .IN8(~na649_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y67     80'h00_0018_00_0040_0A72_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3547_1 ( .OUT(na3547_1), .IN1(1'b1), .IN2(na3356_1), .IN3(na3219_1), .IN4(1'b1), .IN5(na3594_1), .IN6(~na9829_2), .IN7(na8330_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x120y69     80'h00_FE00_00_0000_0CEE_7E00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3548_1 ( .OUT(na3548_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na9940_2), .IN6(na3222_1), .IN7(~na3547_1),
                      .IN8(~na841_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3548_2 ( .OUT(na3548_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3548_1_i) );
// C_MX4a////      x93y100     80'h00_0018_00_0040_0C05_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3549_1 ( .OUT(na3549_1), .IN1(na8332_2), .IN2(1'b0), .IN3(na3276_1), .IN4(1'b0), .IN5(1'b1), .IN6(na3299_2), .IN7(1'b1),
                      .IN8(~na3216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y93     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3550_1 ( .OUT(na3550_1), .IN1(1'b1), .IN2(~na3424_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1434_2), .IN6(na8333_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x108y66     80'h00_0060_00_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3552_4 ( .OUT(na3552_2), .IN1(~na912_1), .IN2(~na450_2), .IN3(~na875_1), .IN4(~na429_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x102y71     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3554_1 ( .OUT(na3554_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na874_1), .IN7(na8339_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3554_2 ( .OUT(na3554_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3554_1_i) );
// C_MX2b////      x117y70     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3555_1 ( .OUT(na3555_1), .IN1(1'b1), .IN2(na3222_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8341_1), .IN8(na841_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x90y80     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3559_1 ( .OUT(na3559_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1598_1), .IN7(1'b1), .IN8(na8346_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a3559_2 ( .OUT(na3559_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3559_1_i) );
// C_///XOR/      x69y86     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3560_4 ( .OUT(na3560_2), .IN1(1'b0), .IN2(na5953_1), .IN3(1'b0), .IN4(na8348_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y77     80'h00_0018_00_0040_0AF1_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3561_1 ( .OUT(na3561_1), .IN1(1'b1), .IN2(~na5953_2), .IN3(1'b1), .IN4(na5955_2), .IN5(~na2389_1), .IN6(na3560_2), .IN7(na10053_2),
                      .IN8(na8349_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x78y86     80'h00_F600_00_0000_0388_73FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a3562_1 ( .OUT(na3562_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na3263_1), .IN7(~na3561_1),
                      .IN8(~na9820_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3562_2 ( .OUT(na3562_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3562_1_i) );
// C_MX4a////      x81y66     80'h00_0018_00_0040_0C4A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3563_1 ( .OUT(na3563_1), .IN1(1'b0), .IN2(na2043_2), .IN3(1'b1), .IN4(na2099_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y62     80'h00_0018_00_0040_0AC2_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3564_1 ( .OUT(na3564_1), .IN1(1'b1), .IN2(na3563_1), .IN3(~na9907_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na1904_2),
                      .IN8(na1987_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y58     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3565_1 ( .OUT(na3565_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5698_2), .IN6(na3564_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x73y78     80'h00_0018_00_0040_0C4A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3566_1 ( .OUT(na3566_1), .IN1(1'b0), .IN2(na2050_2), .IN3(1'b1), .IN4(na2106_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y58     80'h00_0018_00_0040_0AC2_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3567_1 ( .OUT(na3567_1), .IN1(1'b1), .IN2(na3566_1), .IN3(~na9907_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na1922_2),
                      .IN8(na1994_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x71y57     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3568_1 ( .OUT(na3568_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5699_1), .IN6(na3567_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x89y62     80'h00_0018_00_0040_0C4A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3569_1 ( .OUT(na3569_1), .IN1(1'b0), .IN2(na2057_2), .IN3(1'b1), .IN4(na2113_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x73y66     80'h00_0018_00_0040_0AC2_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3570_1 ( .OUT(na3570_1), .IN1(1'b1), .IN2(na3569_1), .IN3(~na9907_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na1932_2),
                      .IN8(na2001_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x73y56     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3571_1 ( .OUT(na3571_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5700_2), .IN6(na3570_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x86y62     80'h00_0018_00_0040_0C4A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3572_1 ( .OUT(na3572_1), .IN1(1'b0), .IN2(na9553_2), .IN3(1'b1), .IN4(na2120_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y70     80'h00_0018_00_0040_0AA1_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3573_1 ( .OUT(na3573_1), .IN1(~na5692_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3572_1), .IN5(1'b1), .IN6(na2008_2), .IN7(1'b0),
                      .IN8(na1942_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x71y56     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3574_1 ( .OUT(na3574_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5701_1), .IN6(na3573_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x82y62     80'h00_0018_00_0040_0C4A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3575_1 ( .OUT(na3575_1), .IN1(1'b0), .IN2(na2071_2), .IN3(1'b1), .IN4(na2127_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y44     80'h00_0018_00_0040_0AA4_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3576_1 ( .OUT(na3576_1), .IN1(~na5692_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3575_1), .IN5(1'b0), .IN6(na1951_2), .IN7(1'b1),
                      .IN8(na2015_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y39     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3577_1 ( .OUT(na3577_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5702_2), .IN6(na3576_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x81y71     80'h00_0018_00_0040_0C4A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3578_1 ( .OUT(na3578_1), .IN1(1'b0), .IN2(na9554_2), .IN3(1'b1), .IN4(na2134_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y46     80'h00_0018_00_0040_0AC2_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3579_1 ( .OUT(na3579_1), .IN1(na3578_1), .IN2(1'b1), .IN3(~na9907_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na9543_2),
                      .IN8(na2022_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y40     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3580_1 ( .OUT(na3580_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5703_1), .IN6(na3579_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x84y67     80'h00_0018_00_0040_0C4A_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3581_1 ( .OUT(na3581_1), .IN1(1'b0), .IN2(na2085_2), .IN3(1'b1), .IN4(na2141_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y48     80'h00_0018_00_0040_0AA4_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3582_1 ( .OUT(na3582_1), .IN1(~na5692_1), .IN2(1'b1), .IN3(na3581_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1969_2), .IN7(1'b1),
                      .IN8(na2029_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y43     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3583_1 ( .OUT(na3583_1), .IN1(na2456_2), .IN2(1'b1), .IN3(1'b1), .IN4(na5705_2), .IN5(na5704_2), .IN6(na3582_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x88y58     80'h00_0018_00_0040_0CEA_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3584_1 ( .OUT(na3584_1), .IN1(1'b0), .IN2(~na2092_2), .IN3(1'b1), .IN4(~na2148_2), .IN5(na5692_1), .IN6(1'b1), .IN7(na5691_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y60     80'h00_0018_00_0040_0AAB_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3585_1 ( .OUT(na3585_1), .IN1(~na5692_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na3584_1), .IN5(1'b1), .IN6(~na2036_2), .IN7(1'b0),
                      .IN8(~na9544_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x87y97     80'h00_0060_00_0000_0C08_FF73
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3586_4 ( .OUT(na3586_2), .IN1(1'b0), .IN2(~na3424_2), .IN3(~na278_1), .IN4(~na3216_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y94     80'h00_0018_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3587_1 ( .OUT(na3587_1), .IN1(~na3354_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3586_2), .IN6(na8352_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//OR/D      x85y87     80'h00_FE00_80_0000_0C8E_3CDA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3588_1 ( .OUT(na3588_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3587_1), .IN7(1'b1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3588_2 ( .OUT(na3588_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3588_1_i) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3588_4 ( .OUT(na3588_2_i), .IN1(na3588_1), .IN2(1'b0), .IN3(~na3550_1), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3588_5 ( .OUT(na3588_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3588_2_i) );
// C_///ORAND/      x115y69     80'h00_0060_00_0000_0C08_FFB7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3589_4 ( .OUT(na3589_2), .IN1(~na3256_1), .IN2(~na3345_1), .IN3(na3218_2), .IN4(~na3590_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x116y74     80'h00_FE00_80_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3590_4 ( .OUT(na3590_2_i), .IN1(~na3589_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3590_5 ( .OUT(na3590_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3590_2_i) );
// C_OR////      x127y116     80'h00_0018_00_0000_0EEE_5A37
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3592_1 ( .OUT(na3592_1), .IN1(~na8357_2), .IN2(~na8152_2), .IN3(1'b0), .IN4(~na8151_1), .IN5(na8357_1), .IN6(1'b0), .IN7(~na8355_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x106y107     80'h00_0060_00_0000_0C0E_FF0B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3593_4 ( .OUT(na3593_2), .IN1(na8358_2), .IN2(~na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x113y67     80'h00_FE00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3594_1 ( .OUT(na3594_1_i), .IN1(1'b1), .IN2(na3343_1), .IN3(1'b1), .IN4(na6626_1), .IN5(na3594_1), .IN6(na9797_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3594_2 ( .OUT(na3594_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3594_1_i) );
// C_MX2b////      x113y69     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3595_1 ( .OUT(na3595_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9822_2), .IN5(~na3352_2), .IN6(1'b0), .IN7(~na3596_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x116y73     80'h00_FE00_80_0000_0C08_FF3D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3596_4 ( .OUT(na3596_2_i), .IN1(~na3595_1), .IN2(na8360_1), .IN3(1'b0), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3596_5 ( .OUT(na3596_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3596_2_i) );
// C_OR////      x75y75     80'h00_0018_00_0000_0CEE_0E00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3597_1 ( .OUT(na3597_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2565_1), .IN6(na8361_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x53y68     80'h00_FA00_80_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3598_4 ( .OUT(na3598_2_i), .IN1(1'b0), .IN2(~na2554_1), .IN3(na2558_1), .IN4(na8363_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3598_5 ( .OUT(na3598_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3598_2_i) );
// C_///ORAND/      x93y97     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3599_4 ( .OUT(na3599_2), .IN1(~na3297_2), .IN2(~na308_1), .IN3(1'b0), .IN4(~na3423_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x95y118     80'h00_FE00_00_0040_0A31_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3600_1 ( .OUT(na3600_1_i), .IN1(~na9823_2), .IN2(1'b1), .IN3(1'b1), .IN4(na6626_1), .IN5(~na3599_2), .IN6(na3600_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3600_2 ( .OUT(na3600_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3600_1_i) );
// C_ORAND////      x76y65     80'h00_0018_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3603_1 ( .OUT(na3603_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na364_2), .IN6(na8370_1), .IN7(na3504_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y88     80'h00_0018_00_0040_0A9C_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3605_1 ( .OUT(na3605_1), .IN1(1'b1), .IN2(~na10054_2), .IN3(1'b1), .IN4(~na9625_2), .IN5(na2570_1), .IN6(1'b0), .IN7(1'b1),
                      .IN8(~na8373_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y80     80'h00_0018_00_0000_0888_C133
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3607_1 ( .OUT(na3607_1), .IN1(1'b1), .IN2(~na8375_2), .IN3(1'b1), .IN4(~na2573_1), .IN5(~na9627_2), .IN6(~na8375_1), .IN7(1'b1),
                      .IN8(na3605_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x76y74     80'h00_0018_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3608_1 ( .OUT(na3608_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na379_1), .IN6(na8377_2), .IN7(~na2558_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x73y65     80'h00_0018_00_0040_0C9C_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3609_1 ( .OUT(na3609_1), .IN1(1'b1), .IN2(1'b0), .IN3(na8378_1), .IN4(~na3608_1), .IN5(1'b1), .IN6(~na3527_1), .IN7(1'b1),
                      .IN8(~na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y84     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3610_4 ( .OUT(na3610_2), .IN1(~na8317_1), .IN2(~na8379_1), .IN3(na1492_1), .IN4(na8319_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x80y66     80'h00_0018_00_0000_0888_FB53
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3611_1 ( .OUT(na3611_1), .IN1(1'b0), .IN2(~na2557_1), .IN3(~na2558_1), .IN4(1'b0), .IN5(na2565_1), .IN6(~na2564_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x80y67     80'h00_0018_00_0040_0C9C_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3612_1 ( .OUT(na3612_1), .IN1(1'b1), .IN2(1'b0), .IN3(na8382_1), .IN4(~na3611_1), .IN5(~na3609_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x121y38     80'h00_0078_00_0020_0C66_A3A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3613_1 ( .OUT(na3613_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na6113_2), .IN7(na9508_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3619_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3613_4 ( .OUT(na3613_2), .COUTY1(na3613_4), .IN1(1'b1), .IN2(~na6113_2), .IN3(na9507_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na6113_2),
                      .IN7(na9508_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3619_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x121y39     80'h00_0078_00_0020_0C66_C3C3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3615_1 ( .OUT(na3615_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na6113_2), .IN7(1'b1), .IN8(na1429_2),
                      .CINX(1'b0), .CINY1(na3613_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3615_4 ( .OUT(na3615_2), .COUTY1(na3615_4), .IN1(1'b1), .IN2(~na6113_2), .IN3(1'b1), .IN4(na1429_1), .IN5(1'b1), .IN6(~na6113_2),
                      .IN7(1'b1), .IN8(na1429_2), .CINX(1'b0), .CINY1(na3613_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x121y40     80'h00_0018_00_0010_0666_003A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3617_1 ( .OUT(na3617_1), .COUTY1(na3617_4), .IN1(na1430_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6117_1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3615_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x122y43     80'h00_0078_00_0020_0C66_ACFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3618_1 ( .OUT(na3618_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na6113_2), .IN7(na9508_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3620_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3618_4 ( .OUT(na3618_2), .COUTY1(na3618_4), .IN1(na1427_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6113_2),
                      .IN7(na9508_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3620_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x121y37     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3619_2 ( .OUT(na3619_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3619_6 ( .COUTY1(na3619_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3619_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x122y42     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3620_2 ( .OUT(na3620_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3620_6 ( .COUTY1(na3620_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3620_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x121y41     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3621_1 ( .OUT(na3621_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3617_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x122y44     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3640_1 ( .OUT(na3640_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1429_2),
                      .CINX(1'b0), .CINY1(na3618_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3640_4 ( .OUT(na3640_2), .COUTY1(na3640_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1429_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1429_2), .CINX(1'b0), .CINY1(na3618_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x122y45     80'h00_0078_00_0020_0C66_5A30
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3644_1 ( .OUT(na3644_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1430_1), .IN6(1'b1), .IN7(~na4072_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3640_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3644_4 ( .OUT(na3644_2), .COUTY1(na3644_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4074_1), .IN5(na1430_1), .IN6(1'b1),
                      .IN7(~na4072_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3640_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x122y46     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3646_1 ( .OUT(na3646_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3644_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x120y37     80'h00_0078_00_0020_0C66_5530
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3651_1 ( .OUT(na3651_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1427_2), .IN6(1'b1), .IN7(~na9507_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3661_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3651_4 ( .OUT(na3651_2), .COUTY1(na3651_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1429_2), .IN5(~na1427_2), .IN6(1'b1),
                      .IN7(~na9507_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3661_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x120y38     80'h00_0078_00_0020_0C66_30F5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3653_1 ( .OUT(na3653_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na1429_1),
                      .CINX(1'b0), .CINY1(na3651_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3653_4 ( .OUT(na3653_2), .COUTY1(na3653_4), .IN1(~na1430_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b1), .IN8(~na1429_1), .CINX(1'b0), .CINY1(na3651_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x134y117     80'h00_0078_00_0020_0C66_3A3A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3655_1 ( .OUT(na3655_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na6055_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na9198_2),
                      .CINX(1'b0), .CINY1(na3662_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3655_4 ( .OUT(na3655_2), .COUTY1(na3655_4), .IN1(na6055_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na9197_2), .IN5(na6055_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(~na9198_2), .CINX(1'b0), .CINY1(na3662_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x134y118     80'h00_0078_00_0020_0C66_5A5A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3657_1 ( .OUT(na3657_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na6055_1), .IN6(1'b1), .IN7(~na320_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3655_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3657_4 ( .OUT(na3657_2), .COUTY1(na3657_4), .IN1(na6055_1), .IN2(1'b1), .IN3(~na320_1), .IN4(1'b1), .IN5(na6055_1), .IN6(1'b1),
                      .IN7(~na320_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3655_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x134y119     80'h00_0018_00_0010_0666_003A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3659_1 ( .OUT(na3659_1), .COUTY1(na3659_4), .IN1(na6055_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na321_2), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3657_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x132y120     80'h00_0078_00_0020_0C66_CAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3660_1 ( .OUT(na3660_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na6055_1), .IN6(1'b1), .IN7(1'b1), .IN8(na9198_2),
                      .CINX(1'b0), .CINY1(na3663_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3660_4 ( .OUT(na3660_2), .COUTY1(na3660_4), .IN1(1'b1), .IN2(na318_1), .IN3(1'b1), .IN4(1'b1), .IN5(na6055_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na9198_2), .CINX(1'b0), .CINY1(na3663_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x120y36     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3661_2 ( .OUT(na3661_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3661_6 ( .COUTY1(na3661_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3661_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x134y116     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3662_2 ( .OUT(na3662_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3662_6 ( .COUTY1(na3662_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3662_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x132y119     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3663_2 ( .OUT(na3663_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3663_6 ( .COUTY1(na3663_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3663_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x120y39     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3664_1 ( .OUT(na3664_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3653_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x134y120     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3665_1 ( .OUT(na3665_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3659_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x132y121     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3682_1 ( .OUT(na3682_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na320_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3660_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3682_4 ( .OUT(na3682_2), .COUTY1(na3682_4), .IN1(1'b1), .IN2(1'b1), .IN3(na320_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na320_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3660_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x132y122     80'h00_0078_00_0020_0C66_C305
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3686_1 ( .OUT(na3686_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na4029_1), .IN7(1'b1), .IN8(na321_2),
                      .CINX(1'b0), .CINY1(na3682_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3686_4 ( .OUT(na3686_2), .COUTY1(na3686_4), .IN1(~na4070_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na4029_1),
                      .IN7(1'b1), .IN8(na321_2), .CINX(1'b0), .CINY1(na3682_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x132y123     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3688_1 ( .OUT(na3688_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3686_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x131y123     80'h00_0078_00_0020_0C66_3350
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3693_1 ( .OUT(na3693_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na318_2), .IN7(1'b1), .IN8(~na9197_2),
                      .CINX(1'b0), .CINY1(na3697_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3693_4 ( .OUT(na3693_2), .COUTY1(na3693_4), .IN1(1'b0), .IN2(1'b0), .IN3(~na320_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na318_2),
                      .IN7(1'b1), .IN8(~na9197_2), .CINX(1'b0), .CINY1(na3697_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x131y124     80'h00_0078_00_0020_0C66_503F
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3695_1 ( .OUT(na3695_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na320_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3693_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3695_4 ( .OUT(na3695_2), .COUTY1(na3695_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na321_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na320_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3693_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x131y122     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3697_2 ( .OUT(na3697_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3697_6 ( .COUTY1(na3697_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3697_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x79y109     80'h00_0078_00_0020_0C66_CAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3698_1 ( .OUT(na3698_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1126_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1864_2),
                      .CINX(1'b0), .CINY1(na3701_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3698_4 ( .OUT(na3698_2), .COUTY1(na3698_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1864_1), .IN5(na1126_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na1864_2), .CINX(1'b0), .CINY1(na3701_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x79y110     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3700_1 ( .OUT(na3700_1), .IN1(na1126_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3698_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x79y108     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3701_2 ( .OUT(na3701_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3701_6 ( .COUTY1(na3701_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3701_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x97y61     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3703_1 ( .OUT(na3703_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1858_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3731_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3703_4 ( .OUT(na3703_2), .COUTY1(na3703_4), .IN1(na456_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1858_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3731_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y62     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3705_1 ( .OUT(na3705_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na464_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3703_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3705_4 ( .OUT(na3705_2), .COUTY1(na3705_4), .IN1(1'b1), .IN2(na470_1), .IN3(1'b0), .IN4(1'b0), .IN5(na464_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3703_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y63     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3707_1 ( .OUT(na3707_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na473_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3705_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3707_4 ( .OUT(na3707_2), .COUTY1(na3707_4), .IN1(na474_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na473_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3705_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y64     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3709_1 ( .OUT(na3709_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na475_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3707_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3709_4 ( .OUT(na3709_2), .COUTY1(na3709_4), .IN1(na476_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na475_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3707_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y65     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3711_1 ( .OUT(na3711_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na477_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3709_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3711_4 ( .OUT(na3711_2), .COUTY1(na3711_4), .IN1(1'b1), .IN2(na1855_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na477_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3709_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y56     80'h00_0078_00_0020_0C66_AAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3712_1 ( .OUT(na3712_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na423_1), .IN6(1'b1), .IN7(na420_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3724_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3712_4 ( .OUT(na3712_2), .COUTY1(na3712_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na424_1), .IN5(na423_1), .IN6(1'b1),
                      .IN7(na420_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3724_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y66     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3714_1 ( .OUT(na3714_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1854_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3711_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3714_4 ( .OUT(na3714_2), .COUTY1(na3714_4), .IN1(na484_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1854_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3711_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y67     80'h00_0078_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3716_1 ( .OUT(na3716_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na485_1),
                      .CINX(1'b0), .CINY1(na3714_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3716_4 ( .OUT(na3716_2), .COUTY1(na3716_4), .IN1(1'b0), .IN2(1'b0), .IN3(na492_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na485_1), .CINX(1'b0), .CINY1(na3714_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y68     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3718_1 ( .OUT(na3718_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na493_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3716_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3718_4 ( .OUT(na3718_2), .COUTY1(na3718_4), .IN1(na494_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na493_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3716_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y69     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3720_1 ( .OUT(na3720_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na495_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3718_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3720_4 ( .OUT(na3720_2), .COUTY1(na3720_4), .IN1(1'b1), .IN2(na496_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na495_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3718_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x97y70     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3722_1 ( .OUT(na3722_1), .COUTY1(na3722_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na497_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na3720_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x97y55     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3724_2 ( .OUT(na3724_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3724_6 ( .COUTY1(na3724_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3724_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x97y57     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3725_1 ( .OUT(na3725_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na437_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3712_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3725_4 ( .OUT(na3725_2), .COUTY1(na3725_4), .IN1(na438_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na437_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3712_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y58     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3727_1 ( .OUT(na3727_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na439_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3725_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3727_4 ( .OUT(na3727_2), .COUTY1(na3727_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na440_1), .IN5(1'b0), .IN6(1'b0), .IN7(na439_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3725_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y59     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3729_1 ( .OUT(na3729_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na441_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3727_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3729_4 ( .OUT(na3729_2), .COUTY1(na3729_4), .IN1(1'b1), .IN2(na442_1), .IN3(1'b0), .IN4(1'b0), .IN5(na441_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3727_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x97y60     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3731_1 ( .OUT(na3731_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na445_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3729_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3731_4 ( .OUT(na3731_2), .COUTY1(na3731_4), .IN1(1'b1), .IN2(na446_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na445_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3729_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x131y125     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3732_1 ( .OUT(na3732_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3695_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x133y101     80'h00_0078_00_0020_0C66_CAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3733_1 ( .OUT(na3733_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na9328_2), .IN6(1'b1), .IN7(1'b1), .IN8(na753_2),
                      .CINX(1'b0), .CINY1(na3740_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3733_4 ( .OUT(na3733_2), .COUTY1(na3733_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na753_1), .IN5(na9328_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na753_2), .CINX(1'b0), .CINY1(na3740_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x133y102     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3735_1 ( .OUT(na3735_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na709_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3733_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3735_4 ( .OUT(na3735_2), .COUTY1(na3735_4), .IN1(1'b0), .IN2(1'b0), .IN3(na709_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na709_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3733_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x133y103     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3737_1 ( .OUT(na3737_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na2953_2),
                      .CINX(1'b0), .CINY1(na3735_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3737_4 ( .OUT(na3737_2), .COUTY1(na3737_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na2953_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na2953_2), .CINX(1'b0), .CINY1(na3735_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x133y104     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3739_1 ( .OUT(na3739_1), .IN1(na2951_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3737_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x133y100     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3740_2 ( .OUT(na3740_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3740_6 ( .COUTY1(na3740_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3740_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x96y115     80'h00_0078_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3742_1 ( .OUT(na3742_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3130_1),
                      .CINX(1'b0), .CINY1(na3771_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3742_4 ( .OUT(na3742_2), .COUTY1(na3742_4), .IN1(1'b1), .IN2(na1656_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na3130_1), .CINX(1'b0), .CINY1(na3771_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y116     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3744_1 ( .OUT(na3744_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3118_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3742_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3744_4 ( .OUT(na3744_2), .COUTY1(na3744_4), .IN1(1'b0), .IN2(1'b0), .IN3(na3113_1), .IN4(1'b1), .IN5(na3118_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3742_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y117     80'h00_0078_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3746_1 ( .OUT(na3746_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3119_1),
                      .CINX(1'b0), .CINY1(na3744_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3746_4 ( .OUT(na3746_2), .COUTY1(na3746_4), .IN1(1'b1), .IN2(na3126_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na3119_1), .CINX(1'b0), .CINY1(na3744_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y118     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3748_1 ( .OUT(na3748_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1695_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3746_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3748_4 ( .OUT(na3748_2), .COUTY1(na3748_4), .IN1(1'b0), .IN2(1'b0), .IN3(na3134_1), .IN4(1'b1), .IN5(na1695_1), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3746_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y119     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3750_1 ( .OUT(na3750_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3139_1),
                      .CINX(1'b0), .CINY1(na3748_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3750_4 ( .OUT(na3750_2), .COUTY1(na3750_4), .IN1(na1903_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na3139_1), .CINX(1'b0), .CINY1(na3748_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y110     80'h00_0078_00_0020_0C66_AAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3751_1 ( .OUT(na3751_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3208_1), .IN6(1'b1), .IN7(na9704_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3772_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3751_4 ( .OUT(na3751_2), .COUTY1(na3751_4), .IN1(1'b0), .IN2(1'b0), .IN3(na3195_1), .IN4(1'b1), .IN5(na3208_1), .IN6(1'b1),
                      .IN7(na9704_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3772_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y120     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3753_1 ( .OUT(na3753_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3147_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3750_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3753_4 ( .OUT(na3753_2), .COUTY1(na3753_4), .IN1(1'b1), .IN2(na3170_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3147_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3750_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y121     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3755_1 ( .OUT(na3755_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3192_1),
                      .CINX(1'b0), .CINY1(na3753_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3755_4 ( .OUT(na3755_2), .COUTY1(na3755_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3201_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na3192_1), .CINX(1'b0), .CINY1(na3753_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y122     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3757_1 ( .OUT(na3757_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3205_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3755_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3757_4 ( .OUT(na3757_2), .COUTY1(na3757_4), .IN1(1'b0), .IN2(1'b0), .IN3(na247_1), .IN4(1'b1), .IN5(1'b1), .IN6(na3205_1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3755_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y123     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3759_1 ( .OUT(na3759_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na2739_1),
                      .CINX(1'b0), .CINY1(na3757_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3759_4 ( .OUT(na3759_2), .COUTY1(na3759_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na322_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na2739_1), .CINX(1'b0), .CINY1(na3757_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y124     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3761_1 ( .OUT(na3761_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2748_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3759_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3761_4 ( .OUT(na3761_2), .COUTY1(na3761_4), .IN1(na2721_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2748_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3759_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x96y125     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3764_1 ( .OUT(na3764_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na2255_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3761_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y111     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3765_1 ( .OUT(na3765_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3190_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3751_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3765_4 ( .OUT(na3765_2), .COUTY1(na3765_4), .IN1(na3169_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3190_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3751_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y112     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3767_1 ( .OUT(na3767_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2157_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3765_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3767_4 ( .OUT(na3767_2), .COUTY1(na3767_4), .IN1(1'b1), .IN2(na3148_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2157_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3765_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y113     80'h00_0078_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3769_1 ( .OUT(na3769_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3146_1),
                      .CINX(1'b0), .CINY1(na3767_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3769_4 ( .OUT(na3769_2), .COUTY1(na3769_4), .IN1(1'b0), .IN2(1'b0), .IN3(na3141_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na3146_1), .CINX(1'b0), .CINY1(na3767_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x96y114     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3771_1 ( .OUT(na3771_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3138_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3769_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3771_4 ( .OUT(na3771_2), .COUTY1(na3771_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1829_1), .IN4(1'b1), .IN5(1'b1), .IN6(na3138_1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3769_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x96y109     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3772_2 ( .OUT(na3772_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3772_6 ( .COUTY1(na3772_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3772_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x127y42     80'h00_0078_00_0020_0C66_0AFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3774_1 ( .OUT(na3774_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3006_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3804_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3774_4 ( .OUT(na3774_2), .COUTY1(na3774_4), .IN1(na3006_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3006_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3804_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y43     80'h00_0078_00_0020_0C66_FC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3776_1 ( .OUT(na3776_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1375_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3774_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3776_4 ( .OUT(na3776_2), .COUTY1(na3776_4), .IN1(1'b1), .IN2(na1375_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1375_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3774_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y44     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3778_1 ( .OUT(na3778_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3003_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3776_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3778_4 ( .OUT(na3778_2), .COUTY1(na3778_4), .IN1(na3003_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3003_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3776_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y45     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3780_1 ( .OUT(na3780_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na1365_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3778_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3780_4 ( .OUT(na3780_2), .COUTY1(na3780_4), .IN1(1'b1), .IN2(1'b1), .IN3(na1365_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1365_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3778_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y46     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3782_1 ( .OUT(na3782_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1260_2),
                      .CINX(1'b0), .CINY1(na3780_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3782_4 ( .OUT(na3782_2), .COUTY1(na3782_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1260_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1260_2), .CINX(1'b0), .CINY1(na3780_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y37     80'h00_0078_00_0020_0C66_CC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3783_1 ( .OUT(na3783_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3026_2), .IN7(1'b1), .IN8(na3027_1),
                      .CINX(1'b0), .CINY1(na3797_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3783_4 ( .OUT(na3783_2), .COUTY1(na3783_4), .IN1(1'b1), .IN2(na3026_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3026_2),
                      .IN7(1'b1), .IN8(na3027_1), .CINX(1'b0), .CINY1(na3797_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y47     80'h00_0078_00_0020_0C66_FC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3785_1 ( .OUT(na3785_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1258_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3782_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3785_4 ( .OUT(na3785_2), .COUTY1(na3785_4), .IN1(1'b1), .IN2(na1258_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1258_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3782_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y48     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3787_1 ( .OUT(na3787_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1256_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3785_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3787_4 ( .OUT(na3787_2), .COUTY1(na3787_4), .IN1(na1256_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1256_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3785_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y49     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3789_1 ( .OUT(na3789_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1254_2),
                      .CINX(1'b0), .CINY1(na3787_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3789_4 ( .OUT(na3789_2), .COUTY1(na3789_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1254_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1254_2), .CINX(1'b0), .CINY1(na3787_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y50     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3791_1 ( .OUT(na3791_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1252_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3789_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3791_4 ( .OUT(na3791_2), .COUTY1(na3791_4), .IN1(na1252_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1252_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3789_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y51     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3793_1 ( .OUT(na3793_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1250_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3791_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3793_4 ( .OUT(na3793_2), .COUTY1(na3793_4), .IN1(1'b1), .IN2(na1250_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1250_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3791_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x127y52     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3796_1 ( .OUT(na3796_1), .COUTY1(na3796_4), .IN1(1'b1), .IN2(na1249_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na3793_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x127y36     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3797_2 ( .OUT(na3797_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3797_6 ( .COUTY1(na3797_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3797_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x127y38     80'h00_0078_00_0020_0C66_AFA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3798_1 ( .OUT(na3798_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3024_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3783_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3798_4 ( .OUT(na3798_2), .COUTY1(na3798_4), .IN1(1'b0), .IN2(1'b0), .IN3(na3024_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3024_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3783_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y39     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3800_1 ( .OUT(na3800_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3022_2),
                      .CINX(1'b0), .CINY1(na3798_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3800_4 ( .OUT(na3800_2), .COUTY1(na3800_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3022_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3022_2), .CINX(1'b0), .CINY1(na3798_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y40     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3802_1 ( .OUT(na3802_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3020_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3800_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3802_4 ( .OUT(na3802_2), .COUTY1(na3802_4), .IN1(1'b1), .IN2(na3020_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3020_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3800_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x127y41     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3804_1 ( .OUT(na3804_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3018_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3802_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3804_4 ( .OUT(na3804_2), .COUTY1(na3804_4), .IN1(1'b1), .IN2(1'b1), .IN3(na3018_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3018_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3802_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x97y71     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3805_1 ( .OUT(na3805_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3722_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y114     80'h00_0078_00_0020_0C66_A0AF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3807_1 ( .OUT(na3807_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3162_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3837_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3807_4 ( .OUT(na3807_2), .COUTY1(na3807_4), .IN1(1'b1), .IN2(1'b1), .IN3(na3162_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3162_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3837_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y115     80'h00_0078_00_0020_0C66_FC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3809_1 ( .OUT(na3809_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3173_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3807_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3809_4 ( .OUT(na3809_2), .COUTY1(na3809_4), .IN1(1'b1), .IN2(na3173_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3173_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3807_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y116     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3811_1 ( .OUT(na3811_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3182_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3809_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3811_4 ( .OUT(na3811_2), .COUTY1(na3811_4), .IN1(na3182_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3182_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3809_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y117     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3813_1 ( .OUT(na3813_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3188_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3811_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3813_4 ( .OUT(na3813_2), .COUTY1(na3813_4), .IN1(1'b1), .IN2(na3188_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3188_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3811_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y118     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3815_1 ( .OUT(na3815_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3115_2),
                      .CINX(1'b0), .CINY1(na3813_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3815_4 ( .OUT(na3815_2), .COUTY1(na3815_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3115_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3115_2), .CINX(1'b0), .CINY1(na3813_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y109     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3816_1 ( .OUT(na3816_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1343_2), .IN7(na3002_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3830_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3816_4 ( .OUT(na3816_2), .COUTY1(na3816_4), .IN1(1'b1), .IN2(na1343_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1343_2),
                      .IN7(na3002_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3830_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y119     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3818_1 ( .OUT(na3818_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3122_2),
                      .CINX(1'b0), .CINY1(na3815_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3818_4 ( .OUT(na3818_2), .COUTY1(na3818_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3122_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3122_2), .CINX(1'b0), .CINY1(na3815_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y120     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3820_1 ( .OUT(na3820_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3127_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3818_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3820_4 ( .OUT(na3820_2), .COUTY1(na3820_4), .IN1(1'b1), .IN2(1'b1), .IN3(na3127_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3127_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3818_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y121     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3822_1 ( .OUT(na3822_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3131_2),
                      .CINX(1'b0), .CINY1(na3820_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3822_4 ( .OUT(na3822_2), .COUTY1(na3822_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3131_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3131_2), .CINX(1'b0), .CINY1(na3820_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y122     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3824_1 ( .OUT(na3824_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3137_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3822_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3824_4 ( .OUT(na3824_2), .COUTY1(na3824_4), .IN1(na3137_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na3137_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3822_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y123     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3826_1 ( .OUT(na3826_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1888_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3824_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3826_4 ( .OUT(na3826_2), .COUTY1(na3826_4), .IN1(1'b1), .IN2(na1888_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1888_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3824_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x48y124     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3829_1 ( .OUT(na3829_1), .COUTY1(na3829_4), .IN1(na3142_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na3826_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x48y108     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3830_2 ( .OUT(na3830_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3830_6 ( .COUTY1(na3830_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3830_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x48y110     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3831_1 ( .OUT(na3831_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2158_2),
                      .CINX(1'b0), .CINY1(na3816_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3831_4 ( .OUT(na3831_2), .COUTY1(na3831_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na2158_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na2158_2), .CINX(1'b0), .CINY1(na3816_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y111     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3833_1 ( .OUT(na3833_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na2692_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3831_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3833_4 ( .OUT(na3833_2), .COUTY1(na3833_4), .IN1(1'b1), .IN2(1'b1), .IN3(na2692_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2692_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3831_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y112     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3835_1 ( .OUT(na3835_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3064_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3833_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3835_4 ( .OUT(na3835_2), .COUTY1(na3835_4), .IN1(1'b1), .IN2(na3064_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3064_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3833_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y113     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3837_1 ( .OUT(na3837_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3159_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3835_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3837_4 ( .OUT(na3837_2), .COUTY1(na3837_4), .IN1(na3159_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3159_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3835_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x127y53     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3838_1 ( .OUT(na3838_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3796_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x111y53     80'h00_0078_00_0020_0C66_AA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3839_1 ( .OUT(na3839_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2996_1), .IN6(1'b1), .IN7(na2995_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3842_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3839_4 ( .OUT(na3839_2), .COUTY1(na3839_4), .IN1(1'b1), .IN2(na2993_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2996_1), .IN6(1'b1),
                      .IN7(na2995_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3842_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x111y54     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3841_1 ( .OUT(na3841_1), .IN1(na2992_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3839_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x111y52     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3842_2 ( .OUT(na3842_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3842_6 ( .COUTY1(na3842_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3842_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x104y54     80'h00_0078_00_0020_0C66_CAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3843_1 ( .OUT(na3843_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1171_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1172_1),
                      .CINX(1'b0), .CINY1(na3846_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3843_4 ( .OUT(na3843_2), .COUTY1(na3843_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1170_1), .IN4(1'b1), .IN5(na1171_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na1172_1), .CINX(1'b0), .CINY1(na3846_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x104y55     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3845_1 ( .OUT(na3845_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1169_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3843_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x104y53     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3846_2 ( .OUT(na3846_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3846_6 ( .COUTY1(na3846_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3846_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x116y44     80'h00_0078_00_0020_0C66_AAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3847_1 ( .OUT(na3847_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1167_1), .IN6(1'b1), .IN7(na1165_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3851_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3847_4 ( .OUT(na3847_2), .COUTY1(na3847_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1165_2), .IN4(1'b1), .IN5(na1167_1), .IN6(1'b1),
                      .IN7(na1165_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3851_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x116y45     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3849_1 ( .OUT(na3849_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1134_2),
                      .CINX(1'b0), .CINY1(na3847_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3849_4 ( .OUT(na3849_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1134_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1134_2),
                      .CINX(1'b0), .CINY1(na3847_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x116y43     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3851_2 ( .OUT(na3851_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3851_6 ( .COUTY1(na3851_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3851_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x82y96     80'h00_0078_00_0020_0C66_AAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3852_1 ( .OUT(na3852_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1187_1), .IN6(1'b1), .IN7(na1186_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3855_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3852_4 ( .OUT(na3852_2), .COUTY1(na3852_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1185_1), .IN4(1'b1), .IN5(na1187_1), .IN6(1'b1),
                      .IN7(na1186_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3855_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x82y97     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3854_1 ( .OUT(na3854_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1184_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3852_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x82y95     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3855_2 ( .OUT(na3855_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3855_6 ( .COUTY1(na3855_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3855_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x84y74     80'h00_0078_00_0020_0C66_AAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3856_1 ( .OUT(na3856_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1222_1), .IN6(1'b1), .IN7(na1221_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3859_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3856_4 ( .OUT(na3856_2), .COUTY1(na3856_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1220_1), .IN4(1'b1), .IN5(na1222_1), .IN6(1'b1),
                      .IN7(na1221_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3859_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x84y75     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3858_1 ( .OUT(na3858_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1219_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3856_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x84y73     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3859_2 ( .OUT(na3859_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3859_6 ( .COUTY1(na3859_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3859_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x82y105     80'h00_0078_00_0020_0C66_AA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3860_1 ( .OUT(na3860_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1193_2), .IN6(1'b1), .IN7(na1191_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3864_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3860_4 ( .OUT(na3860_2), .COUTY1(na3860_4), .IN1(na1193_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1193_2), .IN6(1'b1),
                      .IN7(na1191_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3864_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x82y106     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3862_1 ( .OUT(na3862_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1191_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3860_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3862_4 ( .OUT(na3862_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1188_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1191_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3860_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x82y104     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3864_2 ( .OUT(na3864_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3864_6 ( .COUTY1(na3864_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3864_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x126y103     80'h00_0078_00_0020_0C66_AC0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3865_1 ( .OUT(na3865_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2671_1), .IN7(na2673_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3867_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3865_4 ( .OUT(na3865_2), .IN1(na995_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2671_1), .IN7(na2673_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3867_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x126y102     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3867_2 ( .OUT(na3867_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3867_6 ( .COUTY1(na3867_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3867_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x135y77     80'h00_0078_00_0020_0C66_AAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3868_1 ( .OUT(na3868_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1010_1), .IN6(1'b1), .IN7(na1016_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3870_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3868_4 ( .OUT(na3868_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1018_1), .IN5(na1010_1), .IN6(1'b1), .IN7(na1016_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3870_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x135y76     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3870_2 ( .OUT(na3870_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3870_6 ( .COUTY1(na3870_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3870_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x92y95     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3871_1 ( .OUT(na3871_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na9329_2), .IN6(1'b1), .IN7(1'b1), .IN8(na783_1),
                      .CINX(1'b0), .CINY1(na3873_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3871_4 ( .OUT(na3871_2), .IN1(na2960_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na9329_2), .IN6(1'b1), .IN7(1'b1), .IN8(na783_1),
                      .CINX(1'b0), .CINY1(na3873_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x92y94     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3873_2 ( .OUT(na3873_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3873_6 ( .COUTY1(na3873_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3873_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x133y42     80'h00_0078_00_0020_0C66_AAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3874_1 ( .OUT(na3874_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na790_2), .IN6(1'b1), .IN7(na498_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3877_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3874_4 ( .OUT(na3874_2), .COUTY1(na3874_4), .IN1(1'b0), .IN2(1'b0), .IN3(na498_1), .IN4(1'b1), .IN5(na790_2), .IN6(1'b1),
                      .IN7(na498_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3877_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x133y43     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3876_1 ( .OUT(na3876_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3204_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3874_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x133y41     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3877_2 ( .OUT(na3877_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3877_6 ( .COUTY1(na3877_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3877_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x135y61     80'h00_0078_00_0020_0C66_CAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3878_1 ( .OUT(na3878_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na900_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1333_1),
                      .CINX(1'b0), .CINY1(na3880_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3878_4 ( .OUT(na3878_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1119_1), .IN4(1'b1), .IN5(na900_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1333_1),
                      .CINX(1'b0), .CINY1(na3880_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x135y60     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3880_2 ( .OUT(na3880_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3880_6 ( .COUTY1(na3880_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3880_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x135y45     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3881_1 ( .OUT(na3881_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2718_2), .IN7(na2737_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3884_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3881_4 ( .OUT(na3881_2), .COUTY1(na3881_4), .IN1(1'b1), .IN2(na2718_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2718_2),
                      .IN7(na2737_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3884_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x135y46     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3883_1 ( .OUT(na3883_1), .IN1(na2746_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3881_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x135y44     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3884_2 ( .OUT(na3884_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3884_6 ( .COUTY1(na3884_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3884_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x126y45     80'h00_0078_00_0020_0C66_AAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3885_1 ( .OUT(na3885_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3180_1), .IN6(1'b1), .IN7(na2163_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3887_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3885_4 ( .OUT(na3885_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1727_1), .IN5(na3180_1), .IN6(1'b1), .IN7(na2163_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3887_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x126y44     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3887_2 ( .OUT(na3887_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3887_6 ( .COUTY1(na3887_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3887_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x134y37     80'h00_0078_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3888_1 ( .OUT(na3888_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na985_2), .IN6(1'b1), .IN7(1'b1), .IN8(na9726_2),
                      .CINX(1'b0), .CINY1(na3891_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3888_4 ( .OUT(na3888_2), .COUTY1(na3888_4), .IN1(1'b1), .IN2(na2972_1), .IN3(1'b0), .IN4(1'b0), .IN5(na985_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na9726_2), .CINX(1'b0), .CINY1(na3891_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x134y38     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3890_1 ( .OUT(na3890_1), .IN1(na985_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3888_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x134y36     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3891_2 ( .OUT(na3891_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3891_6 ( .COUTY1(na3891_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3891_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x85y124     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3892_1 ( .OUT(na3892_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na326_2), .IN7(1'b1), .IN8(na1859_2),
                      .CINX(1'b0), .CINY1(na3895_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3892_4 ( .OUT(na3892_2), .COUTY1(na3892_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1859_1), .IN5(1'b1), .IN6(na326_2),
                      .IN7(1'b1), .IN8(na1859_2), .CINX(1'b0), .CINY1(na3895_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x85y125     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3894_1 ( .OUT(na3894_1), .IN1(1'b0), .IN2(1'b0), .IN3(na333_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3892_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x85y123     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3895_2 ( .OUT(na3895_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3895_6 ( .COUTY1(na3895_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3895_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x92y123     80'h00_0078_00_0020_0C66_AA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3896_1 ( .OUT(na3896_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na306_1), .IN6(1'b1), .IN7(na309_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3898_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3896_4 ( .OUT(na3896_2), .IN1(1'b1), .IN2(na311_1), .IN3(1'b0), .IN4(1'b0), .IN5(na306_1), .IN6(1'b1), .IN7(na309_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3898_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x92y122     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3898_2 ( .OUT(na3898_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3898_6 ( .COUTY1(na3898_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3898_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x89y124     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3899_1 ( .OUT(na3899_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na334_1), .IN7(na336_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3902_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3899_4 ( .OUT(na3899_2), .COUTY1(na3899_4), .IN1(1'b0), .IN2(1'b0), .IN3(na336_1), .IN4(1'b1), .IN5(1'b1), .IN6(na334_1),
                      .IN7(na336_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3902_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x89y125     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3901_1 ( .OUT(na3901_1), .IN1(na338_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3899_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x89y123     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3902_2 ( .OUT(na3902_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3902_6 ( .COUTY1(na3902_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3902_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x85y118     80'h00_0078_00_0020_0C66_CAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3903_1 ( .OUT(na3903_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na279_1), .IN6(1'b1), .IN7(1'b1), .IN8(na272_1),
                      .CINX(1'b0), .CINY1(na3905_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3903_4 ( .OUT(na3903_2), .IN1(1'b0), .IN2(1'b0), .IN3(na282_1), .IN4(1'b1), .IN5(na279_1), .IN6(1'b1), .IN7(1'b1), .IN8(na272_1),
                      .CINX(1'b0), .CINY1(na3905_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x85y117     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3905_2 ( .OUT(na3905_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3905_6 ( .COUTY1(na3905_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3905_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x82y123     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3906_1 ( .OUT(na3906_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na291_2), .IN7(na289_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3971_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3906_4 ( .OUT(na3906_2), .COUTY1(na3906_4), .IN1(1'b1), .IN2(na291_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na291_2),
                      .IN7(na289_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3971_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x82y124     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3908_1 ( .OUT(na3908_1), .IN1(1'b0), .IN2(1'b0), .IN3(na289_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3906_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y107     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3909_1 ( .OUT(na3909_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na740_2), .IN6(1'b1), .IN7(1'b1), .IN8(na725_1),
                      .CINX(1'b0), .CINY1(na3974_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3909_4 ( .OUT(na3909_2), .COUTY1(na3909_4), .IN1(na740_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na740_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na725_1), .CINX(1'b0), .CINY1(na3974_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y112     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3910_1 ( .OUT(na3910_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na782_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3937_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3910_4 ( .OUT(na3910_2), .COUTY1(na3910_4), .IN1(1'b0), .IN2(1'b0), .IN3(na782_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na782_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3937_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y113     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3912_1 ( .OUT(na3912_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na795_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3910_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3912_4 ( .OUT(na3912_2), .COUTY1(na3912_4), .IN1(na795_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na795_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3910_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y114     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3914_1 ( .OUT(na3914_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na806_2),
                      .CINX(1'b0), .CINY1(na3912_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3914_4 ( .OUT(na3914_2), .COUTY1(na3914_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na806_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na806_2), .CINX(1'b0), .CINY1(na3912_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y115     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3916_1 ( .OUT(na3916_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na810_2),
                      .CINX(1'b0), .CINY1(na3914_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3916_4 ( .OUT(na3916_2), .COUTY1(na3916_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na810_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na810_2), .CINX(1'b0), .CINY1(na3914_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y116     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3918_1 ( .OUT(na3918_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na822_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3916_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3918_4 ( .OUT(na3918_2), .COUTY1(na3918_4), .IN1(1'b1), .IN2(na822_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na822_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3916_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y117     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3921_1 ( .OUT(na3921_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na826_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3918_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3921_4 ( .OUT(na3921_2), .COUTY1(na3921_4), .IN1(1'b0), .IN2(1'b0), .IN3(na826_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na826_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3918_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y118     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3923_1 ( .OUT(na3923_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na831_2),
                      .CINX(1'b0), .CINY1(na3921_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3923_4 ( .OUT(na3923_2), .COUTY1(na3923_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na831_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na831_2), .CINX(1'b0), .CINY1(na3921_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y119     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3925_1 ( .OUT(na3925_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1497_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3923_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3925_4 ( .OUT(na3925_2), .COUTY1(na3925_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1497_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1497_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3923_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y120     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3927_1 ( .OUT(na3927_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na860_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3925_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3927_4 ( .OUT(na3927_2), .COUTY1(na3927_4), .IN1(na860_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na860_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3925_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y121     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3929_1 ( .OUT(na3929_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na866_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3927_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3929_4 ( .OUT(na3929_2), .IN1(1'b0), .IN2(1'b0), .IN3(na866_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na866_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3927_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y108     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3931_1 ( .OUT(na3931_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na748_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3909_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3931_4 ( .OUT(na3931_2), .COUTY1(na3931_4), .IN1(1'b1), .IN2(na748_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na748_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3909_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y109     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3933_1 ( .OUT(na3933_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1555_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3931_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3933_4 ( .OUT(na3933_2), .COUTY1(na3933_4), .IN1(1'b1), .IN2(na1555_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1555_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3931_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y110     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3935_1 ( .OUT(na3935_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na766_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3933_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3935_4 ( .OUT(na3935_2), .COUTY1(na3935_4), .IN1(na766_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na766_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3933_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x74y111     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3937_1 ( .OUT(na3937_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na774_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3935_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3937_4 ( .OUT(na3937_2), .COUTY1(na3937_4), .IN1(1'b0), .IN2(1'b0), .IN3(na774_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na774_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3935_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x58y55     80'h00_0018_00_0010_0666_00AC
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3939_1 ( .OUT(na3939_1), .COUTY1(na3939_4), .IN1(1'b1), .IN2(na2272_2), .IN3(na2257_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3983_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y63     80'h00_F660_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3941_1 ( .OUT(na3941_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2262_1), .IN7(na2283_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3970_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3941_2 ( .OUT(na3941_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3941_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3941_4 ( .OUT(na3941_2), .COUTY1(na3941_4), .IN1(1'b1), .IN2(na2284_1), .IN3(na2264_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2262_1),
                      .IN7(na2283_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3970_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y64     80'h00_F660_00_0020_0C66_CCAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3943_1 ( .OUT(na3943_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2285_1), .IN7(1'b1), .IN8(na2265_1),
                      .CINX(1'b0), .CINY1(na3941_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3943_2 ( .OUT(na3943_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3943_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3943_4 ( .OUT(na3943_2), .COUTY1(na3943_4), .IN1(na2266_1), .IN2(1'b1), .IN3(na2286_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2285_1),
                      .IN7(1'b1), .IN8(na2265_1), .CINX(1'b0), .CINY1(na3941_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y65     80'h00_F660_00_0020_0C66_AACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3945_1 ( .OUT(na3945_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2267_1), .IN6(1'b1), .IN7(na2287_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3943_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3945_2 ( .OUT(na3945_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3945_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3945_4 ( .OUT(na3945_2), .COUTY1(na3945_4), .IN1(1'b1), .IN2(na2268_1), .IN3(1'b1), .IN4(na2288_1), .IN5(na2267_1), .IN6(1'b1),
                      .IN7(na2287_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3943_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y66     80'h00_F660_00_0020_0C66_AACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3947_1 ( .OUT(na3947_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2269_1), .IN6(1'b1), .IN7(na2289_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3945_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3947_2 ( .OUT(na3947_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3947_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3947_4 ( .OUT(na3947_2), .COUTY1(na3947_4), .IN1(1'b1), .IN2(na2270_1), .IN3(1'b1), .IN4(na2290_1), .IN5(na2269_1), .IN6(1'b1),
                      .IN7(na2289_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3945_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y67     80'h00_F660_00_0020_0C66_CCAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3949_1 ( .OUT(na3949_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2291_1), .IN7(1'b1), .IN8(na2271_1),
                      .CINX(1'b0), .CINY1(na3947_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3949_2 ( .OUT(na3949_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3949_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3949_4 ( .OUT(na3949_2), .COUTY1(na3949_4), .IN1(na5972_1), .IN2(1'b1), .IN3(na2292_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2291_1),
                      .IN7(1'b1), .IN8(na2271_1), .CINX(1'b0), .CINY1(na3947_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF/D///      x58y56     80'h00_F600_00_0010_0666_02A8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3950_1 ( .OUT(na3950_1_i), .COUTY1(na3950_4), .IN1(na9917_2), .IN2(na3263_1), .IN3(na2273_2), .IN4(1'b1), .IN5(na9918_2),
                      .IN6(~na3263_1), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3939_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3950_2 ( .OUT(na3950_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3950_1_i) );
// C_ADDF2/D//ADDF2/      x58y68     80'h00_F660_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3952_1 ( .OUT(na3952_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5972_1), .IN6(1'b1), .IN7(na2293_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3949_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3952_2 ( .OUT(na3952_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3952_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3952_4 ( .OUT(na3952_2), .COUTY1(na3952_4), .IN1(na5972_1), .IN2(1'b1), .IN3(na2294_1), .IN4(1'b1), .IN5(na5972_1), .IN6(1'b1),
                      .IN7(na2293_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3949_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y69     80'h00_F660_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3954_1 ( .OUT(na3954_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5972_1), .IN6(1'b1), .IN7(na2295_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3952_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3954_2 ( .OUT(na3954_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3954_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3954_4 ( .OUT(na3954_2), .COUTY1(na3954_4), .IN1(na5972_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2296_1), .IN5(na5972_1), .IN6(1'b1),
                      .IN7(na2295_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3952_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y70     80'h00_F660_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3956_1 ( .OUT(na3956_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5972_1), .IN6(1'b1), .IN7(na2297_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3954_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3956_2 ( .OUT(na3956_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3956_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3956_4 ( .OUT(na3956_2), .COUTY1(na3956_4), .IN1(na5972_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2298_1), .IN5(na5972_1), .IN6(1'b1),
                      .IN7(na2297_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3954_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y71     80'h00_F660_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3958_1 ( .OUT(na3958_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5972_1), .IN6(1'b1), .IN7(na2299_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3956_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3958_2 ( .OUT(na3958_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3958_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3958_4 ( .OUT(na3958_2), .COUTY1(na3958_4), .IN1(na5972_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2300_1), .IN5(na5972_1), .IN6(1'b1),
                      .IN7(na2299_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3956_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y72     80'h00_F660_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3960_1 ( .OUT(na3960_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5972_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2301_1),
                      .CINX(1'b0), .CINY1(na3958_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3960_2 ( .OUT(na3960_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3960_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3960_4 ( .OUT(na3960_2), .COUTY1(na3960_4), .IN1(na5972_1), .IN2(1'b1), .IN3(na2302_1), .IN4(1'b1), .IN5(na5972_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na2301_1), .CINX(1'b0), .CINY1(na3958_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF/D///      x58y57     80'h00_F600_00_0010_0666_02A8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3961_1 ( .OUT(na3961_1_i), .COUTY1(na3961_4), .IN1(na5963_1), .IN2(na3263_1), .IN3(na2274_1), .IN4(1'b1), .IN5(na5963_2),
                      .IN6(~na3263_1), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3950_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3961_2 ( .OUT(na3961_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3961_1_i) );
// C_ADDF/D///      x58y73     80'h00_F600_00_0010_0666_00AA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3963_1 ( .OUT(na3963_1_i), .IN1(na5972_1), .IN2(1'b1), .IN3(na2303_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3960_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3963_2 ( .OUT(na3963_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3963_1_i) );
// C_ADDF/D///      x58y58     80'h00_F600_00_0010_0666_02A8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3964_1 ( .OUT(na3964_1_i), .COUTY1(na3964_4), .IN1(na9920_2), .IN2(na3263_1), .IN3(na2275_1), .IN4(1'b1), .IN5(na9921_2),
                      .IN6(~na3263_1), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3961_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3964_2 ( .OUT(na3964_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3964_1_i) );
// C_ADDF/D///      x58y59     80'h00_F600_00_0010_0666_02C8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3965_1 ( .OUT(na3965_1_i), .COUTY1(na3965_4), .IN1(na9922_2), .IN2(na3263_1), .IN3(1'b1), .IN4(na2276_1), .IN5(na9923_2),
                      .IN6(~na3263_1), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na3964_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3965_2 ( .OUT(na3965_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3965_1_i) );
// C_ADDF2/D//ADDF2/      x58y60     80'h00_F660_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3966_1 ( .OUT(na3966_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5967_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2277_1),
                      .CINX(1'b0), .CINY1(na3965_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3966_2 ( .OUT(na3966_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3966_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3966_4 ( .OUT(na3966_2), .COUTY1(na3966_4), .IN1(na5967_1), .IN2(1'b1), .IN3(na2278_1), .IN4(1'b1), .IN5(na5967_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na2277_1), .CINX(1'b0), .CINY1(na3965_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y61     80'h00_F660_00_0020_0C66_CACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3968_1 ( .OUT(na3968_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2279_1), .IN6(1'b1), .IN7(1'b1), .IN8(na5969_2),
                      .CINX(1'b0), .CINY1(na3966_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3968_2 ( .OUT(na3968_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3968_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3968_4 ( .OUT(na3968_2), .COUTY1(na3968_4), .IN1(1'b1), .IN2(na2280_1), .IN3(1'b1), .IN4(na5969_1), .IN5(na2279_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na5969_2), .CINX(1'b0), .CINY1(na3966_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x58y62     80'h00_F660_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3970_1 ( .OUT(na3970_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5971_2), .IN6(1'b1), .IN7(na2281_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3968_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3970_2 ( .OUT(na3970_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3970_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3970_4 ( .OUT(na3970_2), .COUTY1(na3970_4), .IN1(na5971_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2282_1), .IN5(na5971_2), .IN6(1'b1),
                      .IN7(na2281_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3968_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x82y122     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3971_2 ( .OUT(na3971_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3971_6 ( .COUTY1(na3971_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3971_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x127y101     80'h00_0078_00_0020_0C66_ACFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3972_1 ( .OUT(na3972_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2671_1), .IN7(na2673_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3988_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3972_4 ( .OUT(na3972_2), .IN1(na995_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2671_1), .IN7(na2673_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3988_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x74y106     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3974_2 ( .OUT(na3974_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3974_6 ( .COUTY1(na3974_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3974_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x134y78     80'h00_0078_00_0020_0C66_AACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3975_1 ( .OUT(na3975_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1010_1), .IN6(1'b1), .IN7(na1016_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4020_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3975_4 ( .OUT(na3975_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1018_1), .IN5(na1010_1), .IN6(1'b1), .IN7(na1016_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4020_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x79y124     80'h00_0078_00_0020_0C66_C5CF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3977_1 ( .OUT(na3977_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3337_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1481_2),
                      .CINX(1'b0), .CINY1(na4025_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3977_4 ( .OUT(na3977_2), .COUTY1(na3977_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1481_1), .IN5(~na3337_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na1481_2), .CINX(1'b0), .CINY1(na4025_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x79y125     80'h00_0018_00_0010_0666_00FA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3979_1 ( .OUT(na3979_1), .IN1(na1392_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3977_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y124     80'h00_0078_00_0020_0C66_A5AF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3980_1 ( .OUT(na3980_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3335_2), .IN6(1'b1), .IN7(na1433_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4026_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3980_4 ( .OUT(na3980_2), .COUTY1(na3980_4), .IN1(1'b1), .IN2(1'b1), .IN3(na1433_1), .IN4(1'b1), .IN5(~na3335_2), .IN6(1'b1),
                      .IN7(na1433_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na4026_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x78y125     80'h00_0018_00_0010_0666_00FC
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a3982_1 ( .OUT(na3982_1), .IN1(1'b1), .IN2(na1414_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3980_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x58y54     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3983_2 ( .OUT(na3983_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3983_6 ( .COUTY1(na3983_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3983_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x45y92     80'h00_FA60_00_0020_0C66_3ACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3984_1 ( .OUT(na3984_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na348_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na2422_1),
                      .CINX(1'b0), .CINY1(na4027_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3984_2 ( .OUT(na3984_1), .CLK(na4116_1), .EN(na347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3984_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3984_4 ( .OUT(na3984_2), .COUTY1(na3984_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na349_1), .IN5(na348_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(~na2422_1), .CINX(1'b0), .CINY1(na4027_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x45y93     80'h00_FA60_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3986_1 ( .OUT(na3986_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na350_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3984_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3986_2 ( .OUT(na3986_1), .CLK(na4116_1), .EN(na347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3986_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3986_4 ( .OUT(na3986_2), .IN1(1'b1), .IN2(na351_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na350_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3984_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x127y100     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3988_2 ( .OUT(na3988_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3988_6 ( .COUTY1(na3988_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3988_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x109y115     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3990_1 ( .OUT(na3990_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1308_1),
                      .CINX(1'b0), .CINY1(na4019_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3990_4 ( .OUT(na3990_2), .COUTY1(na3990_4), .IN1(na1310_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1308_1), .CINX(1'b0), .CINY1(na4019_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y116     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3992_1 ( .OUT(na3992_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1316_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3990_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3992_4 ( .OUT(na3992_2), .COUTY1(na3992_4), .IN1(1'b1), .IN2(na2659_1), .IN3(1'b1), .IN4(1'b1), .IN5(na1316_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3990_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y117     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3994_1 ( .OUT(na3994_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na1318_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3992_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3994_4 ( .OUT(na3994_2), .COUTY1(na3994_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1323_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1318_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na3992_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y118     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3996_1 ( .OUT(na3996_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1325_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3994_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3996_4 ( .OUT(na3996_2), .COUTY1(na3996_4), .IN1(1'b1), .IN2(na1327_1), .IN3(1'b1), .IN4(1'b1), .IN5(na1325_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3994_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y119     80'h00_0078_00_0020_0C66_CFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3998_1 ( .OUT(na3998_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2244_1),
                      .CINX(1'b0), .CINY1(na3996_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3998_4 ( .OUT(na3998_2), .COUTY1(na3998_4), .IN1(1'b1), .IN2(1'b1), .IN3(na2242_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na2244_1), .CINX(1'b0), .CINY1(na3996_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y110     80'h00_0078_00_0020_0C66_CCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a3999_1 ( .OUT(na3999_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1287_1), .IN7(1'b1), .IN8(na1289_1),
                      .CINX(1'b0), .CINY1(na4028_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3999_4 ( .OUT(na3999_2), .COUTY1(na3999_4), .IN1(na1291_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1287_1),
                      .IN7(1'b1), .IN8(na1289_1), .CINX(1'b0), .CINY1(na4028_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y120     80'h00_0078_00_0020_0C66_FCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4001_1 ( .OUT(na4001_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1329_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3998_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4001_4 ( .OUT(na4001_2), .COUTY1(na4001_4), .IN1(na2240_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1329_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3998_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y121     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4003_1 ( .OUT(na4003_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na2237_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4001_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4003_4 ( .OUT(na4003_2), .COUTY1(na4003_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1331_1), .IN5(1'b1), .IN6(1'b1), .IN7(na2237_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4001_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y122     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4005_1 ( .OUT(na4005_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na2235_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4003_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4005_4 ( .OUT(na4005_2), .COUTY1(na4005_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2166_1), .IN5(1'b1), .IN6(1'b1), .IN7(na2235_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4003_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y123     80'h00_0078_00_0020_0C66_FCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4007_1 ( .OUT(na4007_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2161_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4005_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4007_4 ( .OUT(na4007_2), .COUTY1(na4007_4), .IN1(na2159_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2161_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4005_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y124     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4009_1 ( .OUT(na4009_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1335_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4007_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4009_4 ( .OUT(na4009_2), .COUTY1(na4009_4), .IN1(1'b1), .IN2(1'b1), .IN3(na1340_1), .IN4(1'b1), .IN5(na1335_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4007_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x109y125     80'h00_0018_00_0010_0666_00FA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a4012_1 ( .OUT(na4012_1), .IN1(na1901_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na4009_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y111     80'h00_0078_00_0020_0C66_CFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4013_1 ( .OUT(na4013_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1293_1),
                      .CINX(1'b0), .CINY1(na3999_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4013_4 ( .OUT(na4013_2), .COUTY1(na4013_4), .IN1(1'b1), .IN2(1'b1), .IN3(na1295_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1293_1), .CINX(1'b0), .CINY1(na3999_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y112     80'h00_0078_00_0020_0C66_FCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4015_1 ( .OUT(na4015_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1297_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4013_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4015_4 ( .OUT(na4015_2), .COUTY1(na4015_4), .IN1(na1299_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1297_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4013_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y113     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4017_1 ( .OUT(na4017_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1301_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4015_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4017_4 ( .OUT(na4017_2), .COUTY1(na4017_4), .IN1(1'b1), .IN2(1'b1), .IN3(na1303_1), .IN4(1'b1), .IN5(na1301_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4015_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x109y114     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4019_1 ( .OUT(na4019_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2664_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4017_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4019_4 ( .OUT(na4019_2), .COUTY1(na4019_4), .IN1(1'b1), .IN2(1'b1), .IN3(na2662_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2664_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4017_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x134y77     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4020_2 ( .OUT(na4020_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4020_6 ( .COUTY1(na4020_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4020_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x134y123     80'h00_0078_00_0020_0C66_CCA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4021_1 ( .OUT(na4021_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na318_2), .IN7(1'b1), .IN8(na9197_2),
                      .CINX(1'b0), .CINY1(na4030_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4021_4 ( .OUT(na4021_2), .COUTY1(na4021_4), .IN1(1'b0), .IN2(1'b0), .IN3(na320_2), .IN4(1'b1), .IN5(1'b1), .IN6(na318_2),
                      .IN7(1'b1), .IN8(na9197_2), .CINX(1'b0), .CINY1(na4030_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x134y124     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4023_1 ( .OUT(na4023_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na320_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4021_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4023_4 ( .OUT(na4023_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na321_2), .IN5(1'b0), .IN6(1'b0), .IN7(na320_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4021_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x79y123     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4025_2 ( .OUT(na4025_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4025_6 ( .COUTY1(na4025_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4025_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x78y123     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4026_2 ( .OUT(na4026_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4026_6 ( .COUTY1(na4026_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4026_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x45y91     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4027_2 ( .OUT(na4027_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4027_6 ( .COUTY1(na4027_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4027_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x109y109     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4028_2 ( .OUT(na4028_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4028_6 ( .COUTY1(na4028_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4028_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF////      x133y116     80'h00_0018_00_0010_0666_00AA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a4029_1 ( .OUT(na4029_1), .COUTY1(na4029_4), .IN1(na6055_1), .IN2(1'b1), .IN3(na9934_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na4031_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x134y122     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4030_2 ( .OUT(na4030_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4030_6 ( .COUTY1(na4030_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4030_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x133y115     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4031_2 ( .OUT(na4031_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4031_6 ( .COUTY1(na4031_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4031_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x130y86     80'h00_0078_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4033_1 ( .OUT(na4033_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3083_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4062_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4033_4 ( .OUT(na4033_2), .COUTY1(na4033_4), .IN1(na3081_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3083_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4062_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y87     80'h00_0078_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4035_1 ( .OUT(na4035_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3079_1),
                      .CINX(1'b0), .CINY1(na4033_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4035_4 ( .OUT(na4035_2), .COUTY1(na4035_4), .IN1(1'b1), .IN2(na3077_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3079_1), .CINX(1'b0), .CINY1(na4033_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y88     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4037_1 ( .OUT(na4037_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3068_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4035_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4037_4 ( .OUT(na4037_2), .COUTY1(na4037_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1445_1), .IN5(1'b1), .IN6(1'b1), .IN7(na3068_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4035_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y89     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4039_1 ( .OUT(na4039_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3062_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4037_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4039_4 ( .OUT(na4039_2), .COUTY1(na4039_4), .IN1(1'b1), .IN2(na3060_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3062_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4037_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y90     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4041_1 ( .OUT(na4041_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3058_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4039_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4041_4 ( .OUT(na4041_2), .COUTY1(na4041_4), .IN1(1'b1), .IN2(1'b1), .IN3(na3056_1), .IN4(1'b1), .IN5(na3058_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4039_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y81     80'h00_0078_00_0020_0C66_ACCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4042_1 ( .OUT(na4042_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3105_1), .IN7(na3103_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4063_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4042_4 ( .OUT(na4042_2), .COUTY1(na4042_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3101_1), .IN5(1'b1), .IN6(na3105_1),
                      .IN7(na3103_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4063_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y91     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4044_1 ( .OUT(na4044_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3054_1),
                      .CINX(1'b0), .CINY1(na4041_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4044_4 ( .OUT(na4044_2), .COUTY1(na4044_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3052_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3054_1), .CINX(1'b0), .CINY1(na4041_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y92     80'h00_0078_00_0020_0C66_FCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4046_1 ( .OUT(na4046_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3050_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4044_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4046_4 ( .OUT(na4046_2), .COUTY1(na4046_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3048_1), .IN5(1'b1), .IN6(na3050_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4044_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y93     80'h00_0078_00_0020_0C66_FCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4048_1 ( .OUT(na4048_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3046_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4046_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4048_4 ( .OUT(na4048_2), .COUTY1(na4048_4), .IN1(na3044_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3046_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4046_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y94     80'h00_0078_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4050_1 ( .OUT(na4050_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na3042_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4048_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4050_4 ( .OUT(na4050_2), .COUTY1(na4050_4), .IN1(na3040_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3042_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4048_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y95     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4052_1 ( .OUT(na4052_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3038_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4050_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4052_4 ( .OUT(na4052_2), .COUTY1(na4052_4), .IN1(1'b1), .IN2(1'b1), .IN3(na3036_1), .IN4(1'b1), .IN5(1'b1), .IN6(na3038_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4050_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x130y96     80'h00_0018_00_0010_0666_00FA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a4055_1 ( .OUT(na4055_1), .IN1(na3034_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na4052_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y82     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4056_1 ( .OUT(na4056_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3099_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4042_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4056_4 ( .OUT(na4056_2), .COUTY1(na4056_4), .IN1(1'b1), .IN2(1'b1), .IN3(na3097_1), .IN4(1'b1), .IN5(na3099_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4042_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y83     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4058_1 ( .OUT(na4058_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3095_1),
                      .CINX(1'b0), .CINY1(na4056_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4058_4 ( .OUT(na4058_2), .COUTY1(na4058_4), .IN1(na3093_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3095_1), .CINX(1'b0), .CINY1(na4056_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y84     80'h00_0078_00_0020_0C66_FCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4060_1 ( .OUT(na4060_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na3091_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4058_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4060_4 ( .OUT(na4060_2), .COUTY1(na4060_4), .IN1(na3089_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3091_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4058_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x130y85     80'h00_0078_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4062_1 ( .OUT(na4062_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3087_1),
                      .CINX(1'b0), .CINY1(na4060_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4062_4 ( .OUT(na4062_2), .COUTY1(na4062_4), .IN1(1'b1), .IN2(na3085_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na3087_1), .CINX(1'b0), .CINY1(na4060_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x130y80     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4063_2 ( .OUT(na4063_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4063_6 ( .COUTY1(na4063_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4063_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x119y38     80'h00_0078_00_0020_0C66_AAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4064_1 ( .OUT(na4064_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1427_2), .IN6(1'b1), .IN7(na9507_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4068_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4064_4 ( .OUT(na4064_2), .COUTY1(na4064_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1429_2), .IN5(na1427_2), .IN6(1'b1),
                      .IN7(na9507_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na4068_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x119y39     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4066_1 ( .OUT(na4066_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1429_1),
                      .CINX(1'b0), .CINY1(na4064_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4066_4 ( .OUT(na4066_2), .IN1(na1430_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1429_1),
                      .CINX(1'b0), .CINY1(na4064_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x119y37     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4068_2 ( .OUT(na4068_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4068_6 ( .COUTY1(na4068_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4068_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x48y125     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a4069_1 ( .OUT(na4069_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na3829_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x133y117     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a4070_1 ( .OUT(na4070_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na4029_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x124y43     80'h00_0018_00_0010_0666_00CC
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a4072_1 ( .OUT(na4072_1), .COUTY1(na4072_4), .IN1(1'b1), .IN2(na6113_2), .IN3(1'b1), .IN4(na6117_1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na4073_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x124y42     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4073_2 ( .OUT(na4073_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4073_6 ( .COUTY1(na4073_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4073_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x124y44     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a4074_1 ( .OUT(na4074_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na4072_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x125y46     80'h00_0078_00_0020_0C66_CC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4075_1 ( .OUT(na4075_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na9738_2), .IN7(1'b1), .IN8(na3032_2),
                      .CINX(1'b0), .CINY1(na4078_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4075_4 ( .OUT(na4075_2), .COUTY1(na4075_4), .IN1(1'b1), .IN2(na3031_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na9738_2),
                      .IN7(1'b1), .IN8(na3032_2), .CINX(1'b0), .CINY1(na4078_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x125y47     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a4077_1 ( .OUT(na4077_1), .IN1(1'b1), .IN2(na3031_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na4075_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x125y45     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4078_2 ( .OUT(na4078_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4078_6 ( .COUTY1(na4078_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4078_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x132y108     80'h00_0078_00_0020_0C66_AACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4079_1 ( .OUT(na4079_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na8394_1), .IN6(1'b1), .IN7(na10057_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4085_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4079_4 ( .OUT(na4079_2), .COUTY1(na4079_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na8405_1), .IN5(na8394_1), .IN6(1'b1),
                      .IN7(na10057_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na4085_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x132y109     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4081_1 ( .OUT(na4081_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na8405_2),
                      .CINX(1'b0), .CINY1(na4079_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4081_4 ( .OUT(na4081_2), .COUTY1(na4081_4), .IN1(na8416_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na8405_2), .CINX(1'b0), .CINY1(na4079_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x132y110     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4083_1 ( .OUT(na4083_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na8416_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4081_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4083_4 ( .OUT(na4083_2), .IN1(1'b1), .IN2(na8417_1), .IN3(1'b1), .IN4(1'b1), .IN5(na8416_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4081_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x132y107     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4085_2 ( .OUT(na4085_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4085_6 ( .COUTY1(na4085_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4085_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x90y46     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4087_1 ( .OUT(na4087_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2900_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4104_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4087_4 ( .OUT(na4087_2), .COUTY1(na4087_4), .IN1(1'b1), .IN2(na2898_2), .IN3(1'b1), .IN4(1'b1), .IN5(na2900_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4104_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y47     80'h00_0078_00_0020_0C66_CFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4089_1 ( .OUT(na4089_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na301_2),
                      .CINX(1'b0), .CINY1(na4087_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4089_4 ( .OUT(na4089_2), .COUTY1(na4089_4), .IN1(1'b1), .IN2(1'b1), .IN3(na300_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na301_2), .CINX(1'b0), .CINY1(na4087_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y48     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4091_1 ( .OUT(na4091_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na281_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4089_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4091_4 ( .OUT(na4091_2), .COUTY1(na4091_4), .IN1(1'b1), .IN2(na171_1), .IN3(1'b1), .IN4(1'b1), .IN5(na281_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4089_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y49     80'h00_0078_00_0020_0C66_CFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4093_1 ( .OUT(na4093_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2897_1),
                      .CINX(1'b0), .CINY1(na4091_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4093_4 ( .OUT(na4093_2), .COUTY1(na4093_4), .IN1(1'b1), .IN2(1'b1), .IN3(na2899_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na2897_1), .CINX(1'b0), .CINY1(na4091_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x90y50     80'h00_0018_00_0010_0666_00CF
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a4095_1 ( .OUT(na4095_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2897_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na4093_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y41     80'h00_0078_00_0020_0C66_CACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4096_1 ( .OUT(na4096_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2917_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2907_2),
                      .CINX(1'b0), .CINY1(na4105_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4096_4 ( .OUT(na4096_2), .COUTY1(na4096_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2907_1), .IN5(na2917_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na2907_2), .CINX(1'b0), .CINY1(na4105_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y42     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4098_1 ( .OUT(na4098_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na2904_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4096_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4098_4 ( .OUT(na4098_2), .COUTY1(na4098_4), .IN1(1'b1), .IN2(na2904_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2904_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4096_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y43     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4100_1 ( .OUT(na4100_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2901_2),
                      .CINX(1'b0), .CINY1(na4098_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4100_4 ( .OUT(na4100_2), .COUTY1(na4100_4), .IN1(na2902_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na2901_2), .CINX(1'b0), .CINY1(na4098_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y44     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4102_1 ( .OUT(na4102_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2901_1),
                      .CINX(1'b0), .CINY1(na4100_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4102_4 ( .OUT(na4102_2), .COUTY1(na4102_4), .IN1(na2900_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na2901_1), .CINX(1'b0), .CINY1(na4100_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y45     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4104_1 ( .OUT(na4104_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na2899_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4102_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4104_4 ( .OUT(na4104_2), .COUTY1(na4104_4), .IN1(1'b1), .IN2(na2898_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2899_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na4102_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x90y40     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4105_2 ( .OUT(na4105_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4105_6 ( .COUTY1(na4105_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4105_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x117y43     80'h00_0078_00_0020_0C66_AAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4106_1 ( .OUT(na4106_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1167_1), .IN6(1'b1), .IN7(na1165_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4110_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4106_4 ( .OUT(na4106_2), .COUTY1(na4106_4), .IN1(1'b1), .IN2(1'b1), .IN3(na1165_2), .IN4(1'b1), .IN5(na1167_1), .IN6(1'b1),
                      .IN7(na1165_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na4110_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x117y44     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4108_1 ( .OUT(na4108_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2),
                      .CINX(1'b0), .CINY1(na4106_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4108_4 ( .OUT(na4108_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1134_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2),
                      .CINX(1'b0), .CINY1(na4106_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x117y42     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a4110_2 ( .OUT(na4110_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a4110_6 ( .COUTY1(na4110_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na4110_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x83y104     80'h00_0078_00_0020_0C66_AAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4111_1 ( .OUT(na4111_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1193_2), .IN6(1'b1), .IN7(na1191_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na6056_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4111_4 ( .OUT(na4111_2), .COUTY1(na4111_4), .IN1(na1193_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1193_2), .IN6(1'b1),
                      .IN7(na1191_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na6056_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x83y105     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a4113_1 ( .OUT(na4113_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na1191_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4111_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a4113_4 ( .OUT(na4113_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1188_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1191_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na4111_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0000_0014)) 
           _a4116 ( .GLB0(na4116_1), .GLB1(_d0), .GLB2(_d1), .GLB3(_d2), .CLK_FB0(_d3), .CLK_FB1(_d4), .CLK_FB2(_d5), .CLK_FB3(_d6),
                    .CLK0_0(na6627_6), .CLK0_90(na6627_5), .CLK0_180(na6627_4), .CLK0_270(na6627_3), .CLK0_BYP(1'b0), .CLK1_0(1'b0),
                    .CLK1_90(1'b0), .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                    .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                    .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                    .USR_FB3(1'b0) );
// C_AND/DST///      x103y114     80'h20_7500_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4118_1 ( .OUT(na4118_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2725_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0000)) 
           _a4118_2 ( .OUT(na4118_1), .CLK(~na4116_1), .EN(~na3239_1), .SR(~na3_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4118_1_i) );
// C_///AND/DST      x81y37     80'h20_7500_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4119_4 ( .OUT(na4119_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2751_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0100)) 
           _a4119_5 ( .OUT(na4119_2), .CLK(~na4116_1), .EN(~na3275_1), .SR(~na4_2), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4119_2_i) );
// C_AND/D///      x84y57     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4132_1 ( .OUT(na4132_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2996_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4132_2 ( .OUT(na4132_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4132_1_i) );
// C_///AND/D      x82y54     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4133_4 ( .OUT(na4133_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2995_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4133_5 ( .OUT(na4133_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4133_2_i) );
// C_AND/D///      x89y60     80'h00_FE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4134_1 ( .OUT(na4134_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2993_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4134_2 ( .OUT(na4134_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4134_1_i) );
// C_///AND/D      x85y56     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4135_4 ( .OUT(na4135_2_i), .IN1(na2992_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4135_5 ( .OUT(na4135_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4135_2_i) );
// C_AND/D///      x75y74     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4138_1 ( .OUT(na4138_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1187_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4138_2 ( .OUT(na4138_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4138_1_i) );
// C_///AND/D      x79y81     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4139_4 ( .OUT(na4139_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1186_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4139_5 ( .OUT(na4139_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4139_2_i) );
// C_AND/D///      x72y73     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4140_1 ( .OUT(na4140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1185_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4140_2 ( .OUT(na4140_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4140_1_i) );
// C_///AND/D      x80y83     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4141_4 ( .OUT(na4141_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1184_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4141_5 ( .OUT(na4141_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4141_2_i) );
// C_AND/D//AND/D      x133y70     80'h00_FA00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4173_1 ( .OUT(na4173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4173_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4173_2 ( .OUT(na4173_1), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4173_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4173_4 ( .OUT(na4173_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4175_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4173_5 ( .OUT(na4173_2), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4173_2_i) );
// C_AND/D//AND/D      x136y69     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4175_1 ( .OUT(na4175_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4175_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4175_2 ( .OUT(na4175_1), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4175_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4175_4 ( .OUT(na4175_2_i), .IN1(1'b1), .IN2(na4177_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4175_5 ( .OUT(na4175_2), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4175_2_i) );
// C_AND/D//AND/D      x135y68     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4177_1 ( .OUT(na4177_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4177_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4177_2 ( .OUT(na4177_1), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4177_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4177_4 ( .OUT(na4177_2_i), .IN1(1'b1), .IN2(na4179_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4177_5 ( .OUT(na4177_2), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4177_2_i) );
// C_AND/D//AND/D      x131y64     80'h00_FA00_80_0000_0C88_FC5F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4179_1 ( .OUT(na4179_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4179_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4179_2 ( .OUT(na4179_1), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4179_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4179_4 ( .OUT(na4179_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na4204_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4179_5 ( .OUT(na4179_2), .CLK(na4116_1), .EN(na898_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4179_2_i) );
// C_AND/D//AND/D      x120y79     80'h00_FE00_80_0000_0C88_F5AF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4204_1 ( .OUT(na4204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6615_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4204_2 ( .OUT(na4204_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4204_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4204_4 ( .OUT(na4204_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4204_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4204_5 ( .OUT(na4204_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4204_2_i) );
// C_AND/D///      x111y72     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4244_1 ( .OUT(na4244_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na236_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4244_2 ( .OUT(na4244_1), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4244_1_i) );
// C_///AND/D      x114y72     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4245_4 ( .OUT(na4245_2_i), .IN1(1'b1), .IN2(na239_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4245_5 ( .OUT(na4245_2), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4245_2_i) );
// C_AND/D///      x114y72     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4246_1 ( .OUT(na4246_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na240_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4246_2 ( .OUT(na4246_1), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4246_1_i) );
// C_///AND/D      x106y69     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4247_4 ( .OUT(na4247_2_i), .IN1(na241_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4247_5 ( .OUT(na4247_2), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4247_2_i) );
// C_AND/D///      x106y72     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4248_1 ( .OUT(na4248_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na242_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4248_2 ( .OUT(na4248_1), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4248_1_i) );
// C_AND/D///      x108y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4249_1 ( .OUT(na4249_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na243_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4249_2 ( .OUT(na4249_1), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4249_1_i) );
// C_AND/D///      x111y69     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4250_1 ( .OUT(na4250_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na244_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4250_2 ( .OUT(na4250_1), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4250_1_i) );
// C_///AND/D      x113y79     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4251_4 ( .OUT(na4251_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na245_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4251_5 ( .OUT(na4251_2), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4251_2_i) );
// C_AND/D///      x119y81     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4252_1 ( .OUT(na4252_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1013_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4252_2 ( .OUT(na4252_1), .CLK(na4116_1), .EN(na3348_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4252_1_i) );
// C_///AND/D      x111y65     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4253_4 ( .OUT(na4253_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na236_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4253_5 ( .OUT(na4253_2), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4253_2_i) );
// C_AND/D///      x110y69     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4254_1 ( .OUT(na4254_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4254_2 ( .OUT(na4254_1), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4254_1_i) );
// C_///AND/D      x136y47     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4255_4 ( .OUT(na4255_2_i), .IN1(1'b1), .IN2(na240_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4255_5 ( .OUT(na4255_2), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4255_2_i) );
// C_AND/D///      x106y70     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4256_1 ( .OUT(na4256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na241_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4256_2 ( .OUT(na4256_1), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4256_1_i) );
// C_///AND/D      x132y51     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4257_4 ( .OUT(na4257_2_i), .IN1(1'b1), .IN2(na242_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4257_5 ( .OUT(na4257_2), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4257_2_i) );
// C_AND/D///      x130y60     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4258_1 ( .OUT(na4258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na243_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4258_2 ( .OUT(na4258_1), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4258_1_i) );
// C_///AND/D      x123y48     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4259_4 ( .OUT(na4259_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na244_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4259_5 ( .OUT(na4259_2), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4259_2_i) );
// C_///AND/D      x125y44     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4260_4 ( .OUT(na4260_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na245_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4260_5 ( .OUT(na4260_2), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4260_2_i) );
// C_AND/D///      x135y74     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4261_1 ( .OUT(na4261_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1013_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4261_2 ( .OUT(na4261_1), .CLK(na4116_1), .EN(na3350_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4261_1_i) );
// C_///AND/D      x134y47     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4274_4 ( .OUT(na4274_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na236_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4274_5 ( .OUT(na4274_2), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4274_2_i) );
// C_AND/D///      x131y55     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4275_1 ( .OUT(na4275_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na239_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4275_2 ( .OUT(na4275_1), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4275_1_i) );
// C_///AND/D      x131y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4276_4 ( .OUT(na4276_2_i), .IN1(1'b1), .IN2(na240_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4276_5 ( .OUT(na4276_2), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4276_2_i) );
// C_AND/D///      x127y60     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4277_1 ( .OUT(na4277_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na241_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4277_2 ( .OUT(na4277_1), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4277_1_i) );
// C_///AND/D      x135y51     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4278_4 ( .OUT(na4278_2_i), .IN1(1'b1), .IN2(na242_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4278_5 ( .OUT(na4278_2), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4278_2_i) );
// C_///AND/D      x133y54     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4279_4 ( .OUT(na4279_2_i), .IN1(na243_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4279_5 ( .OUT(na4279_2), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4279_2_i) );
// C_///AND/D      x126y48     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4280_4 ( .OUT(na4280_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na244_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4280_5 ( .OUT(na4280_2), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4280_2_i) );
// C_AND/D///      x120y56     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4281_1 ( .OUT(na4281_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na245_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4281_2 ( .OUT(na4281_1), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4281_1_i) );
// C_///AND/D      x134y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4282_4 ( .OUT(na4282_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1013_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4282_5 ( .OUT(na4282_2), .CLK(na4116_1), .EN(na3349_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na4282_2_i) );
// C_AND/D//AND/D      x78y93     80'h00_FE00_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4853_1 ( .OUT(na4853_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6617_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4853_2 ( .OUT(na4853_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4853_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4853_4 ( .OUT(na4853_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4853_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4853_5 ( .OUT(na4853_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4853_2_i) );
// C_AND/D//AND/D      x83y95     80'h00_FE00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4855_1 ( .OUT(na4855_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6604_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4855_2 ( .OUT(na4855_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4855_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4855_4 ( .OUT(na4855_2_i), .IN1(na4855_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4855_5 ( .OUT(na4855_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4855_2_i) );
// C_AND/D///      x116y71     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4856_1 ( .OUT(na4856_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6579_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4856_2 ( .OUT(na4856_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4856_1_i) );
// C_///AND/D      x121y116     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4860_4 ( .OUT(na4860_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na950_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4860_5 ( .OUT(na4860_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4860_2_i) );
// C_AND/D///      x119y74     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4861_1 ( .OUT(na4861_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6580_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4861_2 ( .OUT(na4861_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4861_1_i) );
// C_///AND/D      x117y115     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4864_4 ( .OUT(na4864_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na952_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4864_5 ( .OUT(na4864_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4864_2_i) );
// C_AND/D///      x112y69     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4865_1 ( .OUT(na4865_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6581_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4865_2 ( .OUT(na4865_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4865_1_i) );
// C_///AND/D      x119y116     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4868_4 ( .OUT(na4868_2_i), .IN1(na957_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4868_5 ( .OUT(na4868_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4868_2_i) );
// C_AND/D///      x131y53     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4869_1 ( .OUT(na4869_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6582_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4869_2 ( .OUT(na4869_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4869_1_i) );
// C_///AND/D      x107y116     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4872_4 ( .OUT(na4872_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na959_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4872_5 ( .OUT(na4872_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4872_2_i) );
// C_AND/D///      x136y53     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4873_1 ( .OUT(na4873_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6583_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4873_2 ( .OUT(na4873_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4873_1_i) );
// C_///AND/D      x110y116     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4876_4 ( .OUT(na4876_2_i), .IN1(na970_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4876_5 ( .OUT(na4876_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4876_2_i) );
// C_AND/D//AND/D      x88y114     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4877_1 ( .OUT(na4877_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6572_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4877_2 ( .OUT(na4877_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4877_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4877_4 ( .OUT(na4877_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4877_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4877_5 ( .OUT(na4877_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4877_2_i) );
// C_AND/D///      x131y56     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4878_1 ( .OUT(na4878_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6584_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4878_2 ( .OUT(na4878_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4878_1_i) );
// C_///AND/D      x124y115     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4882_4 ( .OUT(na4882_2_i), .IN1(na968_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4882_5 ( .OUT(na4882_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4882_2_i) );
// C_AND/D///      x132y54     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4883_1 ( .OUT(na4883_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6585_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4883_2 ( .OUT(na4883_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4883_1_i) );
// C_///AND/D      x130y116     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4886_4 ( .OUT(na4886_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na965_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4886_5 ( .OUT(na4886_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4886_2_i) );
// C_AND/D///      x127y55     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4887_1 ( .OUT(na4887_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6586_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4887_2 ( .OUT(na4887_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4887_1_i) );
// C_///AND/D      x113y115     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4890_4 ( .OUT(na4890_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na964_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4890_5 ( .OUT(na4890_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4890_2_i) );
// C_AND/D///      x113y115     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4893_1 ( .OUT(na4893_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na966_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4893_2 ( .OUT(na4893_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4893_1_i) );
// C_AND/D//AND/D      x135y65     80'h00_FE00_80_0000_0C88_FA3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4894_1 ( .OUT(na4894_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6588_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4894_2 ( .OUT(na4894_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4894_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4894_4 ( .OUT(na4894_2_i), .IN1(na4894_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4894_5 ( .OUT(na4894_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4894_2_i) );
// C_AND/D//AND/D      x90y116     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4895_1 ( .OUT(na4895_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6597_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4895_2 ( .OUT(na4895_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4895_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4895_4 ( .OUT(na4895_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4895_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4895_5 ( .OUT(na4895_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4895_2_i) );
// C_AND/D//AND/D      x94y94     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4897_1 ( .OUT(na4897_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6598_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4897_2 ( .OUT(na4897_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4897_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4897_4 ( .OUT(na4897_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4897_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4897_5 ( .OUT(na4897_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4897_2_i) );
// C_AND/D//AND/D      x81y93     80'h00_FE00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4899_1 ( .OUT(na4899_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6569_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4899_2 ( .OUT(na4899_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4899_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4899_4 ( .OUT(na4899_2_i), .IN1(na4899_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4899_5 ( .OUT(na4899_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4899_2_i) );
// C_AND/D//AND/D      x86y110     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4900_1 ( .OUT(na4900_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6599_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4900_2 ( .OUT(na4900_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4900_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4900_4 ( .OUT(na4900_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4900_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4900_5 ( .OUT(na4900_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4900_2_i) );
// C_AND/D//AND/D      x84y114     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4903_1 ( .OUT(na4903_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6600_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4903_2 ( .OUT(na4903_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4903_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4903_4 ( .OUT(na4903_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4903_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4903_5 ( .OUT(na4903_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4903_2_i) );
// C_AND/D//AND/D      x92y116     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4905_1 ( .OUT(na4905_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6601_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4905_2 ( .OUT(na4905_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4905_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4905_4 ( .OUT(na4905_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4905_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4905_5 ( .OUT(na4905_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4905_2_i) );
// C_AND/D//AND/D      x86y112     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4907_1 ( .OUT(na4907_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6602_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4907_2 ( .OUT(na4907_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4907_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4907_4 ( .OUT(na4907_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4907_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4907_5 ( .OUT(na4907_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4907_2_i) );
// C_AND/D//AND/D      x88y84     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4909_1 ( .OUT(na4909_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6593_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4909_2 ( .OUT(na4909_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4909_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4909_4 ( .OUT(na4909_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4909_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4909_5 ( .OUT(na4909_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4909_2_i) );
// C_AND/D//AND/D      x88y82     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4911_1 ( .OUT(na4911_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6594_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4911_2 ( .OUT(na4911_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4911_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4911_4 ( .OUT(na4911_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4911_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4911_5 ( .OUT(na4911_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4911_2_i) );
// C_AND/D//AND/D      x88y88     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4913_1 ( .OUT(na4913_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6595_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4913_2 ( .OUT(na4913_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4913_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4913_4 ( .OUT(na4913_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4913_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4913_5 ( .OUT(na4913_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4913_2_i) );
// C_AND/D//AND/D      x90y90     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4915_1 ( .OUT(na4915_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6596_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4915_2 ( .OUT(na4915_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4915_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4915_4 ( .OUT(na4915_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4915_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4915_5 ( .OUT(na4915_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4915_2_i) );
// C_AND/D//AND/D      x120y74     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4917_1 ( .OUT(na4917_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6574_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4917_2 ( .OUT(na4917_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4917_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4917_4 ( .OUT(na4917_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4917_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4917_5 ( .OUT(na4917_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4917_2_i) );
// C_AND/D//AND/D      x120y72     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4919_1 ( .OUT(na4919_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6575_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4919_2 ( .OUT(na4919_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4919_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4919_4 ( .OUT(na4919_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4919_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4919_5 ( .OUT(na4919_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4919_2_i) );
// C_AND/D//AND/D      x124y78     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4922_1 ( .OUT(na4922_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6573_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4922_2 ( .OUT(na4922_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4922_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4922_4 ( .OUT(na4922_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4922_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4922_5 ( .OUT(na4922_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4922_2_i) );
// C_AND/D//AND/D      x121y117     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4926_1 ( .OUT(na4926_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3333_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4926_2 ( .OUT(na4926_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4926_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4926_4 ( .OUT(na4926_2_i), .IN1(na4926_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4926_5 ( .OUT(na4926_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4926_2_i) );
// C_AND/D//AND/D      x120y113     80'h00_FE00_80_0000_0C88_5FAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4928_1 ( .OUT(na4928_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3333_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4928_2 ( .OUT(na4928_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4928_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4928_4 ( .OUT(na4928_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4928_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4928_5 ( .OUT(na4928_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4928_2_i) );
// C_///AND/D      x122y121     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4930_4 ( .OUT(na4930_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na4928_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4930_5 ( .OUT(na4930_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4930_2_i) );
// C_AND/D///      x123y125     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4933_1 ( .OUT(na4933_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na967_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a4933_2 ( .OUT(na4933_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4933_1_i) );
// C_///AND/D      x115y116     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4936_4 ( .OUT(na4936_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na969_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a4936_5 ( .OUT(na4936_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4936_2_i) );
// C_AND/D///      x115y92     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5167_1 ( .OUT(na5167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3214_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5167_2 ( .OUT(na5167_1), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5167_1_i) );
// C_///AND/D      x109y96     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5168_4 ( .OUT(na5168_2_i), .IN1(na3494_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5168_5 ( .OUT(na5168_2), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5168_2_i) );
// C_AND/D///      x126y109     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5169_1 ( .OUT(na5169_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na107_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5169_2 ( .OUT(na5169_1), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5169_1_i) );
// C_///AND/D      x114y91     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5170_4 ( .OUT(na5170_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na116_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5170_5 ( .OUT(na5170_2), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5170_2_i) );
// C_AND/D///      x121y110     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5171_1 ( .OUT(na5171_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3496_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5171_2 ( .OUT(na5171_1), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5171_1_i) );
// C_///AND/D      x103y96     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5172_4 ( .OUT(na5172_2_i), .IN1(na129_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5172_5 ( .OUT(na5172_2), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5172_2_i) );
// C_AND/D///      x124y116     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5173_1 ( .OUT(na5173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na135_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5173_2 ( .OUT(na5173_1), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5173_1_i) );
// C_///AND/D      x107y95     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5174_4 ( .OUT(na5174_2_i), .IN1(1'b1), .IN2(na142_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5174_5 ( .OUT(na5174_2), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5174_2_i) );
// C_AND/D///      x118y90     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5175_1 ( .OUT(na5175_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na149_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5175_2 ( .OUT(na5175_1), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5175_1_i) );
// C_///AND/D      x119y98     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5176_4 ( .OUT(na5176_2_i), .IN1(na3258_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5176_5 ( .OUT(na5176_2), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5176_2_i) );
// C_AND/D///      x114y99     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5177_1 ( .OUT(na5177_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3499_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5177_2 ( .OUT(na5177_1), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5177_1_i) );
// C_///AND/D      x113y100     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5178_4 ( .OUT(na5178_2_i), .IN1(na103_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5178_5 ( .OUT(na5178_2), .CLK(na4116_1), .EN(na3351_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5178_2_i) );
// C_AND/D//AND/D      x91y114     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5179_1 ( .OUT(na5179_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5179_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5179_2 ( .OUT(na5179_1), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5179_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5179_4 ( .OUT(na5179_2_i), .IN1(1'b1), .IN2(na5181_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5179_5 ( .OUT(na5179_2), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5179_2_i) );
// C_AND/D//AND/D      x93y114     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5181_1 ( .OUT(na5181_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5181_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5181_2 ( .OUT(na5181_1), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5181_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5181_4 ( .OUT(na5181_2_i), .IN1(1'b1), .IN2(na5183_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5181_5 ( .OUT(na5181_2), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5181_2_i) );
// C_AND/D//AND/D      x91y116     80'h00_FA00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5183_1 ( .OUT(na5183_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5183_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5183_2 ( .OUT(na5183_1), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5183_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5183_4 ( .OUT(na5183_2_i), .IN1(na5185_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5183_5 ( .OUT(na5183_2), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5183_2_i) );
// C_AND/D//AND/D      x91y117     80'h00_FA00_80_0000_0C88_FAF3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5185_1 ( .OUT(na5185_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5185_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5185_2 ( .OUT(na5185_1), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5185_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5185_4 ( .OUT(na5185_2_i), .IN1(1'b1), .IN2(~na5223_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5185_5 ( .OUT(na5185_2), .CLK(na4116_1), .EN(na303_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5185_2_i) );
// C_AND/D///      x106y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5215_1 ( .OUT(na5215_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na875_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5215_2 ( .OUT(na5215_1), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5215_1_i) );
// C_///AND/D      x125y54     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5216_4 ( .OUT(na5216_2_i), .IN1(na877_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5216_5 ( .OUT(na5216_2), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5216_2_i) );
// C_AND/D///      x120y61     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5217_1 ( .OUT(na5217_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1894_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5217_2 ( .OUT(na5217_1), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5217_1_i) );
// C_AND/D///      x109y69     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5218_1 ( .OUT(na5218_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1893_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5218_2 ( .OUT(na5218_1), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5218_1_i) );
// C_///AND/D      x129y56     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5219_4 ( .OUT(na5219_2_i), .IN1(na879_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5219_5 ( .OUT(na5219_2), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5219_2_i) );
// C_AND/D///      x117y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5220_1 ( .OUT(na5220_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na880_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5220_2 ( .OUT(na5220_1), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5220_1_i) );
// C_///AND/D      x126y53     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5221_4 ( .OUT(na5221_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na881_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5221_5 ( .OUT(na5221_2), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5221_2_i) );
// C_AND/D///      x118y60     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5222_1 ( .OUT(na5222_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na882_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5222_2 ( .OUT(na5222_1), .CLK(na4116_1), .EN(na3342_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5222_1_i) );
// C_AND/D//AND/D      x91y118     80'h00_FE00_80_0000_0C88_F5FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5223_1 ( .OUT(na5223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6613_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5223_2 ( .OUT(na5223_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5223_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5223_4 ( .OUT(na5223_2_i), .IN1(1'b1), .IN2(na5223_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5223_5 ( .OUT(na5223_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5223_2_i) );
// C_///AND/D      x80y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5228_4 ( .OUT(na5228_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6742_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5228_5 ( .OUT(na5228_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5228_2_i) );
// C_AND/D///      x67y63     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5229_1 ( .OUT(na5229_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6740_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5229_2 ( .OUT(na5229_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5229_1_i) );
// C_///AND/D      x72y68     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5230_4 ( .OUT(na5230_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6739_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5230_5 ( .OUT(na5230_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5230_2_i) );
// C_AND/D///      x68y66     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5231_1 ( .OUT(na5231_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6738_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5231_2 ( .OUT(na5231_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5231_1_i) );
// C_///AND/D      x76y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5232_4 ( .OUT(na5232_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6737_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5232_5 ( .OUT(na5232_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5232_2_i) );
// C_AND/D///      x67y64     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5233_1 ( .OUT(na5233_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6735_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5233_2 ( .OUT(na5233_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5233_1_i) );
// C_///AND/D      x80y63     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5234_4 ( .OUT(na5234_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6734_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5234_5 ( .OUT(na5234_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5234_2_i) );
// C_AND/D///      x67y66     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5235_1 ( .OUT(na5235_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6732_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5235_2 ( .OUT(na5235_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5235_1_i) );
// C_///AND/D      x65y75     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5236_4 ( .OUT(na5236_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6731_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5236_5 ( .OUT(na5236_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5236_2_i) );
// C_AND/D///      x64y73     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5237_1 ( .OUT(na5237_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6730_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5237_2 ( .OUT(na5237_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5237_1_i) );
// C_///AND/D      x64y75     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5238_4 ( .OUT(na5238_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6729_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5238_5 ( .OUT(na5238_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5238_2_i) );
// C_///AND/D      x59y63     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5239_4 ( .OUT(na5239_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6728_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5239_5 ( .OUT(na5239_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5239_2_i) );
// C_AND/D///      x59y65     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5240_1 ( .OUT(na5240_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6726_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5240_2 ( .OUT(na5240_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5240_1_i) );
// C_AND/D///      x68y63     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5241_1 ( .OUT(na5241_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6725_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5241_2 ( .OUT(na5241_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5241_1_i) );
// C_AND/D///      x67y69     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5242_1 ( .OUT(na5242_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6722_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5242_2 ( .OUT(na5242_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5242_1_i) );
// C_///AND/D      x67y69     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5243_4 ( .OUT(na5243_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6721_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5243_5 ( .OUT(na5243_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5243_2_i) );
// C_AND/D///      x57y58     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5244_1 ( .OUT(na5244_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6720_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5244_2 ( .OUT(na5244_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5244_1_i) );
// C_///AND/D      x70y61     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5245_4 ( .OUT(na5245_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6718_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5245_5 ( .OUT(na5245_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5245_2_i) );
// C_AND/D///      x56y67     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5246_1 ( .OUT(na5246_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6717_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5246_2 ( .OUT(na5246_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5246_1_i) );
// C_///AND/D      x65y62     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5247_4 ( .OUT(na5247_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6716_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5247_5 ( .OUT(na5247_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5247_2_i) );
// C_AND/D///      x73y62     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5248_1 ( .OUT(na5248_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6761_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5248_2 ( .OUT(na5248_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5248_1_i) );
// C_///AND/D      x73y57     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5249_4 ( .OUT(na5249_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6760_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5249_5 ( .OUT(na5249_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5249_2_i) );
// C_AND/D///      x67y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5250_1 ( .OUT(na5250_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6758_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5250_2 ( .OUT(na5250_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5250_1_i) );
// C_///AND/D      x73y59     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5251_4 ( .OUT(na5251_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6757_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5251_5 ( .OUT(na5251_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5251_2_i) );
// C_AND/D///      x58y51     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5252_1 ( .OUT(na5252_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6756_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5252_2 ( .OUT(na5252_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5252_1_i) );
// C_///AND/D      x65y55     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5253_4 ( .OUT(na5253_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6755_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5253_5 ( .OUT(na5253_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5253_2_i) );
// C_///AND/D      x68y59     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5254_4 ( .OUT(na5254_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6754_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5254_5 ( .OUT(na5254_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5254_2_i) );
// C_///AND/D      x68y61     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5255_4 ( .OUT(na5255_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6751_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5255_5 ( .OUT(na5255_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5255_2_i) );
// C_AND/D///      x62y53     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5256_1 ( .OUT(na5256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6748_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5256_2 ( .OUT(na5256_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5256_1_i) );
// C_///AND/D      x78y59     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5257_4 ( .OUT(na5257_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6747_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5257_5 ( .OUT(na5257_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5257_2_i) );
// C_AND/D///      x61y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5258_1 ( .OUT(na5258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6746_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5258_2 ( .OUT(na5258_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5258_1_i) );
// C_///AND/D      x75y59     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5259_4 ( .OUT(na5259_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6744_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5259_5 ( .OUT(na5259_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5259_2_i) );
// C_AND/D//AND/D      x73y97     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5261_1 ( .OUT(na5261_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3323_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5261_2 ( .OUT(na5261_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5261_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5261_4 ( .OUT(na5261_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3321_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5261_5 ( .OUT(na5261_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5261_2_i) );
// C_AND/D///      x62y57     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5263_1 ( .OUT(na5263_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6874_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5263_2 ( .OUT(na5263_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5263_1_i) );
// C_///AND/D      x66y53     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5264_4 ( .OUT(na5264_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6873_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5264_5 ( .OUT(na5264_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5264_2_i) );
// C_AND/D///      x66y56     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5265_1 ( .OUT(na5265_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6872_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5265_2 ( .OUT(na5265_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5265_1_i) );
// C_///AND/D      x59y54     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5266_4 ( .OUT(na5266_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6865_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5266_5 ( .OUT(na5266_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5266_2_i) );
// C_AND/D///      x66y62     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5267_1 ( .OUT(na5267_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6863_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5267_2 ( .OUT(na5267_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5267_1_i) );
// C_///AND/D      x57y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5268_4 ( .OUT(na5268_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6862_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5268_5 ( .OUT(na5268_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5268_2_i) );
// C_AND/D///      x61y62     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5269_1 ( .OUT(na5269_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6861_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5269_2 ( .OUT(na5269_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5269_1_i) );
// C_///AND/D      x61y62     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5270_4 ( .OUT(na5270_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6860_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5270_5 ( .OUT(na5270_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5270_2_i) );
// C_AND/D///      x56y56     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5271_1 ( .OUT(na5271_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6858_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5271_2 ( .OUT(na5271_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5271_1_i) );
// C_///AND/D      x59y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5272_4 ( .OUT(na5272_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6857_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5272_5 ( .OUT(na5272_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5272_2_i) );
// C_///AND/D      x55y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5273_4 ( .OUT(na5273_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6856_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5273_5 ( .OUT(na5273_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5273_2_i) );
// C_///AND/D      x67y56     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5274_4 ( .OUT(na5274_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6854_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5274_5 ( .OUT(na5274_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5274_2_i) );
// C_AND/D///      x57y60     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5275_1 ( .OUT(na5275_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6852_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5275_2 ( .OUT(na5275_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5275_1_i) );
// C_///AND/D      x59y58     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5276_4 ( .OUT(na5276_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6851_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5276_5 ( .OUT(na5276_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5276_2_i) );
// C_AND/D///      x59y60     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5277_1 ( .OUT(na5277_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6850_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5277_2 ( .OUT(na5277_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5277_1_i) );
// C_///AND/D      x55y58     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5278_4 ( .OUT(na5278_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6848_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5278_5 ( .OUT(na5278_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5278_2_i) );
// C_AND/D///      x57y62     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5279_1 ( .OUT(na5279_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6846_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5279_2 ( .OUT(na5279_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5279_1_i) );
// C_AND/D///      x65y62     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5280_1 ( .OUT(na5280_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6844_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5280_2 ( .OUT(na5280_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5280_1_i) );
// C_///AND/D      x57y60     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5281_4 ( .OUT(na5281_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6843_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5281_5 ( .OUT(na5281_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5281_2_i) );
// C_///AND/D      x59y64     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5282_4 ( .OUT(na5282_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6842_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5282_5 ( .OUT(na5282_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5282_2_i) );
// C_AND/D///      x59y58     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5283_1 ( .OUT(na5283_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6895_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5283_2 ( .OUT(na5283_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5283_1_i) );
// C_AND/D///      x67y56     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5284_1 ( .OUT(na5284_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6894_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5284_2 ( .OUT(na5284_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5284_1_i) );
// C_///AND/D      x65y56     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5285_4 ( .OUT(na5285_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6893_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5285_5 ( .OUT(na5285_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5285_2_i) );
// C_AND/D///      x68y58     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5286_1 ( .OUT(na5286_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6890_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5286_2 ( .OUT(na5286_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5286_1_i) );
// C_AND/D///      x68y56     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5287_1 ( .OUT(na5287_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6885_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5287_2 ( .OUT(na5287_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5287_1_i) );
// C_///AND/D      x55y44     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5288_4 ( .OUT(na5288_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6884_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5288_5 ( .OUT(na5288_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5288_2_i) );
// C_///AND/D      x61y52     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5289_4 ( .OUT(na5289_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5289_5 ( .OUT(na5289_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5289_2_i) );
// C_///AND/D      x55y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5290_4 ( .OUT(na5290_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6882_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5290_5 ( .OUT(na5290_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5290_2_i) );
// C_AND/D///      x55y50     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5291_1 ( .OUT(na5291_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6880_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5291_2 ( .OUT(na5291_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5291_1_i) );
// C_///AND/D      x61y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5292_4 ( .OUT(na5292_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6878_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5292_5 ( .OUT(na5292_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5292_2_i) );
// C_AND/D///      x57y50     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5293_1 ( .OUT(na5293_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6877_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5293_2 ( .OUT(na5293_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5293_1_i) );
// C_///AND/D      x53y48     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5294_4 ( .OUT(na5294_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6876_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5294_5 ( .OUT(na5294_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5294_2_i) );
// C_AND/D///      x77y70     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5402_1 ( .OUT(na5402_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5953_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5402_2 ( .OUT(na5402_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5402_1_i) );
// C_///AND/D      x76y74     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5403_4 ( .OUT(na5403_2_i), .IN1(1'b1), .IN2(na5953_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5403_5 ( .OUT(na5403_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5403_2_i) );
// C_AND/D//AND/D      x68y112     80'h00_FE00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5435_1 ( .OUT(na5435_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5261_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5435_2 ( .OUT(na5435_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5435_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5435_4 ( .OUT(na5435_2_i), .IN1(na5261_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5435_5 ( .OUT(na5435_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5435_2_i) );
// C_AND/D///      x93y94     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5445_1 ( .OUT(na5445_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na568_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5445_2 ( .OUT(na5445_1), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5445_1_i) );
// C_///AND/D      x100y103     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5446_4 ( .OUT(na5446_2_i), .IN1(na1897_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5446_5 ( .OUT(na5446_2), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5446_2_i) );
// C_AND/D///      x89y110     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5447_1 ( .OUT(na5447_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na894_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5447_2 ( .OUT(na5447_1), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5447_1_i) );
// C_///AND/D      x102y95     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5448_4 ( .OUT(na5448_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na897_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5448_5 ( .OUT(na5448_2), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5448_2_i) );
// C_AND/D///      x90y112     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5449_1 ( .OUT(na5449_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na902_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5449_2 ( .OUT(na5449_1), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5449_1_i) );
// C_AND/D///      x88y110     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5450_1 ( .OUT(na5450_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1364_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5450_2 ( .OUT(na5450_1), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5450_1_i) );
// C_///AND/D      x97y91     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5451_4 ( .OUT(na5451_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1366_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5451_5 ( .OUT(na5451_2), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5451_2_i) );
// C_AND/D///      x87y112     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5452_1 ( .OUT(na5452_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na895_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5452_2 ( .OUT(na5452_1), .CLK(na4116_1), .EN(na3353_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5452_1_i) );
// C_AND/D///      x74y101     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5456_1 ( .OUT(na5456_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6498_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5456_2 ( .OUT(na5456_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5456_1_i) );
// C_AND/D///      x76y97     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5457_1 ( .OUT(na5457_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6499_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5457_2 ( .OUT(na5457_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5457_1_i) );
// C_///AND/D      x72y99     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5458_4 ( .OUT(na5458_2_i), .IN1(na6500_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5458_5 ( .OUT(na5458_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5458_2_i) );
// C_AND/D///      x75y100     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5459_1 ( .OUT(na5459_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6501_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5459_2 ( .OUT(na5459_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5459_1_i) );
// C_AND/D///      x70y101     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5460_1 ( .OUT(na5460_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6502_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5460_2 ( .OUT(na5460_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5460_1_i) );
// C_///AND/D      x76y97     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5461_4 ( .OUT(na5461_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6503_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5461_5 ( .OUT(na5461_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5461_2_i) );
// C_///AND/D      x70y83     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5462_4 ( .OUT(na5462_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6504_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5462_5 ( .OUT(na5462_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5462_2_i) );
// C_AND/D///      x80y97     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5463_1 ( .OUT(na5463_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6505_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5463_2 ( .OUT(na5463_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5463_1_i) );
// C_AND/D///      x72y101     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5464_1 ( .OUT(na5464_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6506_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5464_2 ( .OUT(na5464_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5464_1_i) );
// C_AND/D///      x78y97     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5465_1 ( .OUT(na5465_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6507_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5465_2 ( .OUT(na5465_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5465_1_i) );
// C_///AND/D      x72y101     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5466_4 ( .OUT(na5466_2_i), .IN1(na6508_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5466_5 ( .OUT(na5466_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5466_2_i) );
// C_///AND/D      x79y98     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5467_4 ( .OUT(na5467_2_i), .IN1(na6509_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5467_5 ( .OUT(na5467_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5467_2_i) );
// C_AND/D///      x68y109     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5468_1 ( .OUT(na5468_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6510_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5468_2 ( .OUT(na5468_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5468_1_i) );
// C_AND/D///      x66y107     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5469_1 ( .OUT(na5469_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6511_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5469_2 ( .OUT(na5469_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5469_1_i) );
// C_///AND/D      x70y105     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5470_4 ( .OUT(na5470_2_i), .IN1(1'b1), .IN2(na6512_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5470_5 ( .OUT(na5470_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5470_2_i) );
// C_AND/D///      x70y95     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5471_1 ( .OUT(na5471_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6513_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5471_2 ( .OUT(na5471_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5471_1_i) );
// C_///AND/D      x70y101     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5472_4 ( .OUT(na5472_2_i), .IN1(1'b1), .IN2(na6514_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5472_5 ( .OUT(na5472_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5472_2_i) );
// C_AND/D///      x58y97     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5473_1 ( .OUT(na5473_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6515_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5473_2 ( .OUT(na5473_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5473_1_i) );
// C_///AND/D      x68y105     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5474_4 ( .OUT(na5474_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6516_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5474_5 ( .OUT(na5474_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5474_2_i) );
// C_AND/D///      x66y99     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5475_1 ( .OUT(na5475_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6517_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5475_2 ( .OUT(na5475_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5475_1_i) );
// C_///AND/D      x70y107     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5476_4 ( .OUT(na5476_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6518_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5476_5 ( .OUT(na5476_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5476_2_i) );
// C_AND/D///      x68y105     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5477_1 ( .OUT(na5477_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6519_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5477_2 ( .OUT(na5477_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5477_1_i) );
// C_///AND/D      x76y101     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5478_4 ( .OUT(na5478_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6520_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5478_5 ( .OUT(na5478_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5478_2_i) );
// C_AND/D///      x66y105     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5479_1 ( .OUT(na5479_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6521_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5479_2 ( .OUT(na5479_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5479_1_i) );
// C_///AND/D      x72y105     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5480_4 ( .OUT(na5480_2_i), .IN1(1'b1), .IN2(na6522_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5480_5 ( .OUT(na5480_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5480_2_i) );
// C_AND/D///      x70y105     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5481_1 ( .OUT(na5481_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6523_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5481_2 ( .OUT(na5481_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5481_1_i) );
// C_///AND/D      x74y101     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5482_4 ( .OUT(na5482_2_i), .IN1(1'b1), .IN2(na6524_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5482_5 ( .OUT(na5482_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5482_2_i) );
// C_AND/D///      x68y107     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5483_1 ( .OUT(na5483_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6525_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5483_2 ( .OUT(na5483_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5483_1_i) );
// C_///AND/D      x76y105     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5484_4 ( .OUT(na5484_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5484_5 ( .OUT(na5484_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5484_2_i) );
// C_AND/D///      x72y105     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5485_1 ( .OUT(na5485_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6527_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5485_2 ( .OUT(na5485_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5485_1_i) );
// C_///AND/D      x84y97     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5486_4 ( .OUT(na5486_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6528_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5486_5 ( .OUT(na5486_2), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5486_2_i) );
// C_AND/D///      x72y103     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5487_1 ( .OUT(na5487_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6529_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5487_2 ( .OUT(na5487_1), .CLK(na4116_1), .EN(na404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5487_1_i) );
// C_///AND/D      x50y92     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5488_4 ( .OUT(na5488_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6308_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5488_5 ( .OUT(na5488_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5488_2_i) );
// C_AND/D///      x59y78     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5489_1 ( .OUT(na5489_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6309_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5489_2 ( .OUT(na5489_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5489_1_i) );
// C_///AND/D      x55y82     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5490_4 ( .OUT(na5490_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6310_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5490_5 ( .OUT(na5490_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5490_2_i) );
// C_AND/D///      x55y81     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5491_1 ( .OUT(na5491_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6324_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5491_2 ( .OUT(na5491_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5491_1_i) );
// C_///AND/D      x56y83     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5492_4 ( .OUT(na5492_2_i), .IN1(na6312_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5492_5 ( .OUT(na5492_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5492_2_i) );
// C_///AND/D      x54y86     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5493_4 ( .OUT(na5493_2_i), .IN1(na6313_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5493_5 ( .OUT(na5493_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5493_2_i) );
// C_///AND/D      x47y91     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5494_4 ( .OUT(na5494_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6314_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5494_5 ( .OUT(na5494_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5494_2_i) );
// C_AND/D///      x53y81     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5495_1 ( .OUT(na5495_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6315_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5495_2 ( .OUT(na5495_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5495_1_i) );
// C_///AND/D      x48y92     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5496_4 ( .OUT(na5496_2_i), .IN1(na6325_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5496_5 ( .OUT(na5496_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5496_2_i) );
// C_AND/D///      x56y83     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5497_1 ( .OUT(na5497_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6317_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5497_2 ( .OUT(na5497_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5497_1_i) );
// C_///AND/D      x47y95     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5498_4 ( .OUT(na5498_2_i), .IN1(na6318_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5498_5 ( .OUT(na5498_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5498_2_i) );
// C_AND/D///      x47y90     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5499_1 ( .OUT(na5499_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6319_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5499_2 ( .OUT(na5499_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5499_1_i) );
// C_///AND/D      x50y95     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5500_4 ( .OUT(na5500_2_i), .IN1(na6320_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5500_5 ( .OUT(na5500_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5500_2_i) );
// C_AND/D///      x48y90     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5501_1 ( .OUT(na5501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6321_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5501_2 ( .OUT(na5501_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5501_1_i) );
// C_///AND/D      x49y89     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5502_4 ( .OUT(na5502_2_i), .IN1(na6322_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5502_5 ( .OUT(na5502_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5502_2_i) );
// C_AND/D///      x49y91     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5503_1 ( .OUT(na5503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6323_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5503_2 ( .OUT(na5503_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5503_1_i) );
// C_///AND/D      x45y88     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5504_4 ( .OUT(na5504_2_i), .IN1(na6324_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5504_5 ( .OUT(na5504_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5504_2_i) );
// C_AND/D///      x48y91     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5505_1 ( .OUT(na5505_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6325_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5505_2 ( .OUT(na5505_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5505_1_i) );
// C_///AND/D      x49y91     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5506_4 ( .OUT(na5506_2_i), .IN1(na6326_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5506_5 ( .OUT(na5506_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5506_2_i) );
// C_AND/D///      x49y90     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5507_1 ( .OUT(na5507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6327_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5507_2 ( .OUT(na5507_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5507_1_i) );
// C_///AND/D      x57y98     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5508_4 ( .OUT(na5508_2_i), .IN1(na6328_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5508_5 ( .OUT(na5508_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5508_2_i) );
// C_AND/D///      x48y94     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5509_1 ( .OUT(na5509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6329_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5509_2 ( .OUT(na5509_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5509_1_i) );
// C_///AND/D      x51y94     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5510_4 ( .OUT(na5510_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6330_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5510_5 ( .OUT(na5510_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5510_2_i) );
// C_AND/D///      x49y93     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5511_1 ( .OUT(na5511_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6331_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5511_2 ( .OUT(na5511_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5511_1_i) );
// C_///AND/D      x62y101     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5512_4 ( .OUT(na5512_2_i), .IN1(na6332_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5512_5 ( .OUT(na5512_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5512_2_i) );
// C_AND/D///      x48y96     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5513_1 ( .OUT(na5513_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6333_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5513_2 ( .OUT(na5513_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5513_1_i) );
// C_///AND/D      x49y93     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5514_4 ( .OUT(na5514_2_i), .IN1(na6334_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5514_5 ( .OUT(na5514_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5514_2_i) );
// C_AND/D///      x50y95     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5515_1 ( .OUT(na5515_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6335_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5515_2 ( .OUT(na5515_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5515_1_i) );
// C_///AND/D      x67y83     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5516_4 ( .OUT(na5516_2_i), .IN1(na6336_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5516_5 ( .OUT(na5516_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5516_2_i) );
// C_AND/D///      x50y96     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5517_1 ( .OUT(na5517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6320_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5517_2 ( .OUT(na5517_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5517_1_i) );
// C_///AND/D      x63y108     80'h00_F600_80_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5518_4 ( .OUT(na5518_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na404_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5518_5 ( .OUT(na5518_2), .CLK(na4116_1), .EN(~na359_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5518_2_i) );
// C_AND/D///      x82y72     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5585_1 ( .OUT(na5585_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5946_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5585_2 ( .OUT(na5585_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5585_1_i) );
// C_///AND/D      x79y70     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5586_4 ( .OUT(na5586_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5228_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5586_5 ( .OUT(na5586_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5586_2_i) );
// C_AND/D///      x78y68     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5587_1 ( .OUT(na5587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5229_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5587_2 ( .OUT(na5587_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5587_1_i) );
// C_///AND/D      x83y66     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5588_4 ( .OUT(na5588_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5230_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5588_5 ( .OUT(na5588_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5588_2_i) );
// C_AND/D///      x78y67     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5589_1 ( .OUT(na5589_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5231_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5589_2 ( .OUT(na5589_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5589_1_i) );
// C_///AND/D      x73y60     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5590_4 ( .OUT(na5590_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5232_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5590_5 ( .OUT(na5590_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5590_2_i) );
// C_AND/D///      x75y61     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5591_1 ( .OUT(na5591_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5233_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5591_2 ( .OUT(na5591_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5591_1_i) );
// C_///AND/D      x71y62     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5592_4 ( .OUT(na5592_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5234_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5592_5 ( .OUT(na5592_2), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5592_2_i) );
// C_AND/D///      x73y58     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5593_1 ( .OUT(na5593_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5235_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5593_2 ( .OUT(na5593_1), .CLK(na4116_1), .EN(~na523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5593_1_i) );
// C_AND/D//AND/D      x52y37     80'h00_FE00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5684_1 ( .OUT(na5684_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5684_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5684_2 ( .OUT(na5684_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5684_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5684_4 ( .OUT(na5684_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5931_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5684_5 ( .OUT(na5684_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5684_2_i) );
// C_AND/D//AND/D      x52y40     80'h00_FE00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5685_1 ( .OUT(na5685_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5685_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5685_2 ( .OUT(na5685_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5685_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5685_4 ( .OUT(na5685_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5932_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5685_5 ( .OUT(na5685_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5685_2_i) );
// C_AND/D//AND/D      x51y37     80'h00_FE00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5686_1 ( .OUT(na5686_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5686_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5686_2 ( .OUT(na5686_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5686_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5686_4 ( .OUT(na5686_2_i), .IN1(na5935_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5686_5 ( .OUT(na5686_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5686_2_i) );
// C_AND/D//AND/D      x53y36     80'h00_FE00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5687_1 ( .OUT(na5687_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5687_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5687_2 ( .OUT(na5687_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5687_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5687_4 ( .OUT(na5687_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5932_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5687_5 ( .OUT(na5687_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5687_2_i) );
// C_AND/D//AND/D      x50y35     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5688_1 ( .OUT(na5688_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5688_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5688_2 ( .OUT(na5688_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5688_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5688_4 ( .OUT(na5688_2_i), .IN1(na5935_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5688_5 ( .OUT(na5688_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5688_2_i) );
// C_///AND/D      x81y46     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5689_4 ( .OUT(na5689_2_i), .IN1(na356_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5689_5 ( .OUT(na5689_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5689_2_i) );
// C_AND/D///      x77y72     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5690_1 ( .OUT(na5690_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na354_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5690_2 ( .OUT(na5690_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5690_1_i) );
// C_AND/D//AND/D      x86y41     80'h00_FE00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5691_1 ( .OUT(na5691_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5689_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5691_2 ( .OUT(na5691_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5691_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5691_4 ( .OUT(na5691_2_i), .IN1(na5936_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5691_5 ( .OUT(na5691_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5691_2_i) );
// C_AND/D//AND/D      x85y41     80'h00_FE00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5692_1 ( .OUT(na5692_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5690_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5692_2 ( .OUT(na5692_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5692_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5692_4 ( .OUT(na5692_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5692_5 ( .OUT(na5692_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5692_2_i) );
// C_///AND/D      x50y86     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5695_4 ( .OUT(na5695_2_i), .IN1(1'b1), .IN2(na3984_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5695_5 ( .OUT(na5695_2), .CLK(na4116_1), .EN(na347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5695_2_i) );
// C_AND/D///      x50y87     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5697_1 ( .OUT(na5697_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3986_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5697_2 ( .OUT(na5697_1), .CLK(na4116_1), .EN(na347_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5697_1_i) );
// C_///AND/D      x71y67     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5698_4 ( .OUT(na5698_2_i), .IN1(1'b1), .IN2(na2594_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5698_5 ( .OUT(na5698_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5698_2_i) );
// C_AND/D///      x73y67     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5699_1 ( .OUT(na5699_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2596_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5699_2 ( .OUT(na5699_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5699_1_i) );
// C_///AND/D      x73y67     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5700_4 ( .OUT(na5700_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2597_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5700_5 ( .OUT(na5700_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5700_2_i) );
// C_AND/D///      x73y71     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5701_1 ( .OUT(na5701_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2598_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5701_2 ( .OUT(na5701_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5701_1_i) );
// C_///AND/D      x73y71     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5702_4 ( .OUT(na5702_2_i), .IN1(na2599_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5702_5 ( .OUT(na5702_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5702_2_i) );
// C_AND/D///      x71y67     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5703_1 ( .OUT(na5703_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2600_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5703_2 ( .OUT(na5703_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5703_1_i) );
// C_///AND/D      x71y69     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5704_4 ( .OUT(na5704_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2601_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5704_5 ( .OUT(na5704_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5704_2_i) );
// C_AND/D//AND/D      x62y42     80'h00_FE00_80_0000_0C88_CF5F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5705_1 ( .OUT(na5705_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2602_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5705_2 ( .OUT(na5705_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5705_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5705_4 ( .OUT(na5705_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na403_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5705_5 ( .OUT(na5705_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5705_2_i) );
// C_AND/D///      x63y66     80'h00_FE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5706_1 ( .OUT(na5706_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2603_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5706_2 ( .OUT(na5706_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5706_1_i) );
// C_///AND/D      x68y69     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5707_4 ( .OUT(na5707_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2604_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5707_5 ( .OUT(na5707_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5707_2_i) );
// C_///AND/D      x73y75     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5708_4 ( .OUT(na5708_2_i), .IN1(na2605_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5708_5 ( .OUT(na5708_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5708_2_i) );
// C_///AND/D      x65y69     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5709_4 ( .OUT(na5709_2_i), .IN1(na2606_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5709_5 ( .OUT(na5709_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5709_2_i) );
// C_AND/D///      x70y73     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5710_1 ( .OUT(na5710_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2607_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5710_2 ( .OUT(na5710_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5710_1_i) );
// C_///AND/D      x69y76     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5711_4 ( .OUT(na5711_2_i), .IN1(1'b1), .IN2(na2608_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5711_5 ( .OUT(na5711_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5711_2_i) );
// C_///AND/D      x74y77     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5712_4 ( .OUT(na5712_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2609_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5712_5 ( .OUT(na5712_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5712_2_i) );
// C_AND/D///      x71y69     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5713_1 ( .OUT(na5713_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2610_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5713_2 ( .OUT(na5713_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5713_1_i) );
// C_///AND/D      x71y68     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5714_4 ( .OUT(na5714_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2611_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5714_5 ( .OUT(na5714_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5714_2_i) );
// C_AND/D///      x67y74     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5715_1 ( .OUT(na5715_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2612_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5715_2 ( .OUT(na5715_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5715_1_i) );
// C_///AND/D      x75y74     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5716_4 ( .OUT(na5716_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2613_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5716_5 ( .OUT(na5716_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5716_2_i) );
// C_///AND/D      x65y76     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5717_4 ( .OUT(na5717_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2614_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5717_5 ( .OUT(na5717_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5717_2_i) );
// C_///AND/D      x73y72     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5718_4 ( .OUT(na5718_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2615_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5718_5 ( .OUT(na5718_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5718_2_i) );
// C_///AND/D      x71y70     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5719_4 ( .OUT(na5719_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2616_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5719_5 ( .OUT(na5719_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5719_2_i) );
// C_///AND/D      x73y70     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5720_4 ( .OUT(na5720_2_i), .IN1(1'b1), .IN2(na2617_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5720_5 ( .OUT(na5720_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5720_2_i) );
// C_AND/D///      x67y78     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5721_1 ( .OUT(na5721_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2618_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5721_2 ( .OUT(na5721_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5721_1_i) );
// C_AND/D///      x71y74     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5722_1 ( .OUT(na5722_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2619_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5722_2 ( .OUT(na5722_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5722_1_i) );
// C_AND/D///      x69y76     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5723_1 ( .OUT(na5723_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2620_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5723_2 ( .OUT(na5723_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5723_1_i) );
// C_///AND/D      x69y74     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5724_4 ( .OUT(na5724_2_i), .IN1(1'b1), .IN2(na2621_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5724_5 ( .OUT(na5724_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5724_2_i) );
// C_AND/D///      x63y78     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5725_1 ( .OUT(na5725_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2622_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5725_2 ( .OUT(na5725_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5725_1_i) );
// C_///AND/D      x79y78     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5726_4 ( .OUT(na5726_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2623_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5726_5 ( .OUT(na5726_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5726_2_i) );
// C_///AND/D      x77y80     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5727_4 ( .OUT(na5727_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2624_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5727_5 ( .OUT(na5727_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5727_2_i) );
// C_AND/D///      x71y72     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5728_1 ( .OUT(na5728_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2625_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5728_2 ( .OUT(na5728_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5728_1_i) );
// C_AND/D///      x71y70     80'h00_FE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5729_1 ( .OUT(na5729_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2626_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5729_2 ( .OUT(na5729_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5729_1_i) );
// C_///AND/D      x71y102     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5795_4 ( .OUT(na5795_2_i), .IN1(na740_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5795_5 ( .OUT(na5795_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5795_2_i) );
// C_AND/D///      x71y102     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5796_1 ( .OUT(na5796_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na740_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5796_2 ( .OUT(na5796_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5796_1_i) );
// C_///AND/D      x68y102     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5797_4 ( .OUT(na5797_2_i), .IN1(1'b1), .IN2(na748_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5797_5 ( .OUT(na5797_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5797_2_i) );
// C_///AND/D      x69y92     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5798_4 ( .OUT(na5798_2_i), .IN1(1'b1), .IN2(na748_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5798_5 ( .OUT(na5798_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5798_2_i) );
// C_AND/D///      x55y97     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5799_1 ( .OUT(na5799_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1555_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5799_2 ( .OUT(na5799_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5799_1_i) );
// C_///AND/D      x56y97     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5800_4 ( .OUT(na5800_2_i), .IN1(1'b1), .IN2(na1555_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5800_5 ( .OUT(na5800_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5800_2_i) );
// C_AND/D///      x54y97     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5801_1 ( .OUT(na5801_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na766_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5801_2 ( .OUT(na5801_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5801_1_i) );
// C_///AND/D      x55y98     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5802_4 ( .OUT(na5802_2_i), .IN1(na766_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5802_5 ( .OUT(na5802_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5802_2_i) );
// C_AND/D///      x56y97     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5803_1 ( .OUT(na5803_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na774_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5803_2 ( .OUT(na5803_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5803_1_i) );
// C_///AND/D      x71y95     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5804_4 ( .OUT(na5804_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na774_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5804_5 ( .OUT(na5804_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5804_2_i) );
// C_///AND/D      x54y97     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5805_4 ( .OUT(na5805_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na782_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5805_5 ( .OUT(na5805_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5805_2_i) );
// C_///AND/D      x55y97     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5806_4 ( .OUT(na5806_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na782_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5806_5 ( .OUT(na5806_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5806_2_i) );
// C_AND/D///      x55y98     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5807_1 ( .OUT(na5807_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na795_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5807_2 ( .OUT(na5807_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5807_1_i) );
// C_AND/D///      x59y98     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5808_1 ( .OUT(na5808_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na795_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5808_2 ( .OUT(na5808_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5808_1_i) );
// C_///AND/D      x72y94     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5809_4 ( .OUT(na5809_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na806_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5809_5 ( .OUT(na5809_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5809_2_i) );
// C_AND/D///      x54y99     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5810_1 ( .OUT(na5810_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na806_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5810_2 ( .OUT(na5810_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5810_1_i) );
// C_///AND/D      x68y97     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5811_4 ( .OUT(na5811_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na810_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5811_5 ( .OUT(na5811_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5811_2_i) );
// C_///AND/D      x66y103     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5812_4 ( .OUT(na5812_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na810_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5812_5 ( .OUT(na5812_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5812_2_i) );
// C_///AND/D      x71y104     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5813_4 ( .OUT(na5813_2_i), .IN1(1'b1), .IN2(na822_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5813_5 ( .OUT(na5813_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5813_2_i) );
// C_AND/D///      x66y104     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5814_1 ( .OUT(na5814_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na822_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5814_2 ( .OUT(na5814_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5814_1_i) );
// C_///AND/D      x74y105     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5815_4 ( .OUT(na5815_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na826_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5815_5 ( .OUT(na5815_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5815_2_i) );
// C_AND/D///      x62y91     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5816_1 ( .OUT(na5816_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na826_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5816_2 ( .OUT(na5816_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5816_1_i) );
// C_///AND/D      x62y91     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5817_4 ( .OUT(na5817_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na831_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5817_5 ( .OUT(na5817_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5817_2_i) );
// C_///AND/D      x67y95     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5818_4 ( .OUT(na5818_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na831_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5818_5 ( .OUT(na5818_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5818_2_i) );
// C_AND/D///      x66y109     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5819_1 ( .OUT(na5819_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1497_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5819_2 ( .OUT(na5819_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5819_1_i) );
// C_///AND/D      x54y99     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5820_4 ( .OUT(na5820_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1497_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5820_5 ( .OUT(na5820_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5820_2_i) );
// C_AND/D///      x58y100     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5821_1 ( .OUT(na5821_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na860_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5821_2 ( .OUT(na5821_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5821_1_i) );
// C_///AND/D      x62y94     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5822_4 ( .OUT(na5822_2_i), .IN1(na860_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5822_5 ( .OUT(na5822_2), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5822_2_i) );
// C_AND/D///      x62y94     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5823_1 ( .OUT(na5823_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na866_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5823_2 ( .OUT(na5823_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5823_1_i) );
// C_AND/D///      x57y100     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5824_1 ( .OUT(na5824_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na866_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5824_2 ( .OUT(na5824_1), .CLK(na4116_1), .EN(~na343_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5824_1_i) );
// C_///AND/D      x71y89     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5830_4 ( .OUT(na5830_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3966_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5830_5 ( .OUT(na5830_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5830_2_i) );
// C_AND/D///      x67y79     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5832_1 ( .OUT(na5832_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3968_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5832_2 ( .OUT(na5832_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5832_1_i) );
// C_AND/D///      x73y84     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5834_1 ( .OUT(na5834_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3970_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5834_2 ( .OUT(na5834_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5834_1_i) );
// C_///AND/D      x74y89     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5836_4 ( .OUT(na5836_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3941_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5836_5 ( .OUT(na5836_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5836_2_i) );
// C_AND/D///      x74y87     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5838_1 ( .OUT(na5838_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3943_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5838_2 ( .OUT(na5838_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5838_1_i) );
// C_AND/D///      x74y83     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5840_1 ( .OUT(na5840_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3945_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5840_2 ( .OUT(na5840_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5840_1_i) );
// C_AND/D///      x74y85     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5842_1 ( .OUT(na5842_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3947_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5842_2 ( .OUT(na5842_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5842_1_i) );
// C_///AND/D      x72y91     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5844_4 ( .OUT(na5844_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3949_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5844_5 ( .OUT(na5844_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5844_2_i) );
// C_///AND/D      x73y85     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5846_4 ( .OUT(na5846_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3952_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5846_5 ( .OUT(na5846_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5846_2_i) );
// C_AND/D///      x73y90     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5848_1 ( .OUT(na5848_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3954_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5848_2 ( .OUT(na5848_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5848_1_i) );
// C_///AND/D      x75y91     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5850_4 ( .OUT(na5850_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3956_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5850_5 ( .OUT(na5850_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5850_2_i) );
// C_AND/D///      x74y89     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5852_1 ( .OUT(na5852_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3958_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5852_2 ( .OUT(na5852_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5852_1_i) );
// C_AND/D///      x75y92     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5854_1 ( .OUT(na5854_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3960_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5854_2 ( .OUT(na5854_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5854_1_i) );
// C_///AND/D      x52y100     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5888_4 ( .OUT(na5888_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5488_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5888_5 ( .OUT(na5888_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5888_2_i) );
// C_AND/D///      x56y99     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5889_1 ( .OUT(na5889_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5489_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5889_2 ( .OUT(na5889_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5889_1_i) );
// C_///AND/D      x52y98     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5890_4 ( .OUT(na5890_2_i), .IN1(1'b1), .IN2(na5490_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5890_5 ( .OUT(na5890_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5890_2_i) );
// C_AND/D///      x48y100     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5891_1 ( .OUT(na5891_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5491_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5891_2 ( .OUT(na5891_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5891_1_i) );
// C_///AND/D      x48y100     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5892_4 ( .OUT(na5892_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5492_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5892_5 ( .OUT(na5892_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5892_2_i) );
// C_AND/D///      x46y103     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5893_1 ( .OUT(na5893_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5493_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5893_2 ( .OUT(na5893_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5893_1_i) );
// C_///AND/D      x46y100     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5894_4 ( .OUT(na5894_2_i), .IN1(na5494_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5894_5 ( .OUT(na5894_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5894_2_i) );
// C_AND/D///      x46y98     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5895_1 ( .OUT(na5895_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5495_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5895_2 ( .OUT(na5895_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5895_1_i) );
// C_///AND/D      x44y100     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5896_4 ( .OUT(na5896_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5496_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5896_5 ( .OUT(na5896_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5896_2_i) );
// C_AND/D///      x47y100     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5897_1 ( .OUT(na5897_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5497_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5897_2 ( .OUT(na5897_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5897_1_i) );
// C_///AND/D      x46y104     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5898_4 ( .OUT(na5898_2_i), .IN1(na5498_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5898_5 ( .OUT(na5898_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5898_2_i) );
// C_AND/D///      x48y98     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5899_1 ( .OUT(na5899_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5499_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5899_2 ( .OUT(na5899_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5899_1_i) );
// C_///AND/D      x50y108     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5900_4 ( .OUT(na5900_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5500_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5900_5 ( .OUT(na5900_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5900_2_i) );
// C_AND/D///      x44y98     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5901_1 ( .OUT(na5901_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5501_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5901_2 ( .OUT(na5901_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5901_1_i) );
// C_///AND/D      x48y98     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5902_4 ( .OUT(na5902_2_i), .IN1(na5502_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5902_5 ( .OUT(na5902_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5902_2_i) );
// C_AND/D///      x50y100     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5903_1 ( .OUT(na5903_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5503_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5903_2 ( .OUT(na5903_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5903_1_i) );
// C_///AND/D      x46y98     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5904_4 ( .OUT(na5904_2_i), .IN1(1'b1), .IN2(na5504_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5904_5 ( .OUT(na5904_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5904_2_i) );
// C_AND/D///      x46y100     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5905_1 ( .OUT(na5905_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5505_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5905_2 ( .OUT(na5905_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5905_1_i) );
// C_///AND/D      x50y98     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5906_4 ( .OUT(na5906_2_i), .IN1(na5506_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5906_5 ( .OUT(na5906_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5906_2_i) );
// C_AND/D///      x52y98     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5907_1 ( .OUT(na5907_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5507_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5907_2 ( .OUT(na5907_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5907_1_i) );
// C_///AND/D      x56y98     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5908_4 ( .OUT(na5908_2_i), .IN1(1'b1), .IN2(na5508_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5908_5 ( .OUT(na5908_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5908_2_i) );
// C_AND/D///      x50y98     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5909_1 ( .OUT(na5909_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5509_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5909_2 ( .OUT(na5909_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5909_1_i) );
// C_///AND/D      x50y100     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5910_4 ( .OUT(na5910_2_i), .IN1(1'b1), .IN2(na5510_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5910_5 ( .OUT(na5910_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5910_2_i) );
// C_AND/D///      x52y100     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5911_1 ( .OUT(na5911_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5511_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5911_2 ( .OUT(na5911_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5911_1_i) );
// C_///AND/D      x56y120     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5912_4 ( .OUT(na5912_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5512_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5912_5 ( .OUT(na5912_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5912_2_i) );
// C_AND/D///      x46y102     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5913_1 ( .OUT(na5913_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5513_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5913_2 ( .OUT(na5913_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5913_1_i) );
// C_///AND/D      x48y102     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5914_4 ( .OUT(na5914_2_i), .IN1(na5514_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5914_5 ( .OUT(na5914_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5914_2_i) );
// C_AND/D///      x50y102     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5915_1 ( .OUT(na5915_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5515_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5915_2 ( .OUT(na5915_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5915_1_i) );
// C_///AND/D      x56y100     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5916_4 ( .OUT(na5916_2_i), .IN1(na5516_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5916_5 ( .OUT(na5916_2), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5916_2_i) );
// C_AND/D///      x44y100     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5917_1 ( .OUT(na5917_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5517_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5917_2 ( .OUT(na5917_1), .CLK(na4116_1), .EN(~na404_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5917_1_i) );
// C_///AND/D      x68y71     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5925_4 ( .OUT(na5925_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5938_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5925_5 ( .OUT(na5925_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5925_2_i) );
// C_///AND/D      x54y101     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5926_4 ( .OUT(na5926_2_i), .IN1(1'b1), .IN2(na5939_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5926_5 ( .OUT(na5926_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5926_2_i) );
// C_AND/D///      x53y99     80'h00_FE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5927_1 ( .OUT(na5927_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5940_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5927_2 ( .OUT(na5927_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5927_1_i) );
// C_AND/D///      x79y85     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5930_1 ( .OUT(na5930_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5946_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5930_2 ( .OUT(na5930_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5930_1_i) );
// C_///AND/D      x76y50     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5931_4 ( .OUT(na5931_2_i), .IN1(1'b1), .IN2(na5948_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5931_5 ( .OUT(na5931_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5931_2_i) );
// C_AND/D//AND/D      x56y45     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5932_1 ( .OUT(na5932_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5962_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5932_2 ( .OUT(na5932_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5932_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5932_4 ( .OUT(na5932_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5964_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5932_5 ( .OUT(na5932_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5932_2_i) );
// C_AND/D//AND/D      x55y43     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5935_1 ( .OUT(na5935_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5965_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5935_2 ( .OUT(na5935_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5935_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5935_4 ( .OUT(na5935_2_i), .IN1(na5963_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5935_5 ( .OUT(na5935_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5935_2_i) );
// C_AND/D///      x79y73     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5936_1 ( .OUT(na5936_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5953_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5936_2 ( .OUT(na5936_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5936_1_i) );
// C_///AND/D      x86y57     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5937_4 ( .OUT(na5937_2_i), .IN1(1'b1), .IN2(na5953_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5937_5 ( .OUT(na5937_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5937_2_i) );
// C_AND/D///      x76y50     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5938_1 ( .OUT(na5938_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5955_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5938_2 ( .OUT(na5938_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5938_1_i) );
// C_///AND/D      x73y88     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5939_4 ( .OUT(na5939_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5969_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5939_5 ( .OUT(na5939_2), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5939_2_i) );
// C_AND/D///      x69y86     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5940_1 ( .OUT(na5940_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5971_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5940_2 ( .OUT(na5940_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5940_1_i) );
// C_///AND/D      x88y68     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5941_4 ( .OUT(na5941_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2552_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5941_5 ( .OUT(na5941_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5941_2_i) );
// C_AND/D///      x77y67     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5942_1 ( .OUT(na5942_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2553_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5942_2 ( .OUT(na5942_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5942_1_i) );
// C_///AND/D      x77y83     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5943_4 ( .OUT(na5943_2_i), .IN1(1'b1), .IN2(na2554_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5943_5 ( .OUT(na5943_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5943_2_i) );
// C_AND/D///      x73y69     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5944_1 ( .OUT(na5944_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2555_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5944_2 ( .OUT(na5944_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5944_1_i) );
// C_///AND/D      x80y85     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5945_4 ( .OUT(na5945_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5945_5 ( .OUT(na5945_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5945_2_i) );
// C_AND/D///      x81y73     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5946_1 ( .OUT(na5946_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2557_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5946_2 ( .OUT(na5946_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5946_1_i) );
// C_///AND/D      x78y88     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5947_4 ( .OUT(na5947_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2558_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5947_5 ( .OUT(na5947_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5947_2_i) );
// C_AND/D///      x65y56     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5948_1 ( .OUT(na5948_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2559_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5948_2 ( .OUT(na5948_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5948_1_i) );
// C_AND/D//AND/D      x71y94     80'h00_FA00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5953_1 ( .OUT(na5953_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2564_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5953_2 ( .OUT(na5953_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5953_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5953_4 ( .OUT(na5953_2_i), .IN1(na2565_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5953_5 ( .OUT(na5953_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5953_2_i) );
// C_///AND/D      x74y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5955_4 ( .OUT(na5955_2_i), .IN1(na2566_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5955_5 ( .OUT(na5955_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5955_2_i) );
// C_AND/D///      x55y64     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5956_1 ( .OUT(na5956_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2574_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5956_2 ( .OUT(na5956_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5956_1_i) );
// C_///AND/D      x67y66     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5957_4 ( .OUT(na5957_2_i), .IN1(na2576_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5957_5 ( .OUT(na5957_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5957_2_i) );
// C_AND/D///      x53y65     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5958_1 ( .OUT(na5958_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2578_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5958_2 ( .OUT(na5958_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5958_1_i) );
// C_///AND/D      x61y68     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5959_4 ( .OUT(na5959_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2580_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5959_5 ( .OUT(na5959_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5959_2_i) );
// C_AND/D///      x53y68     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5960_1 ( .OUT(na5960_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2582_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5960_2 ( .OUT(na5960_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5960_1_i) );
// C_///AND/D      x70y76     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5961_4 ( .OUT(na5961_2_i), .IN1(na2584_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5961_5 ( .OUT(na5961_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5961_2_i) );
// C_AND/D//AND/D      x62y60     80'h00_FA00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5962_1 ( .OUT(na5962_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5962_2 ( .OUT(na5962_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5962_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5962_4 ( .OUT(na5962_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2560_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5962_5 ( .OUT(na5962_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5962_2_i) );
// C_AND/D//AND/D      x63y59     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5963_1 ( .OUT(na5963_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2588_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5963_2 ( .OUT(na5963_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5963_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5963_4 ( .OUT(na5963_2_i), .IN1(1'b1), .IN2(na2561_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5963_5 ( .OUT(na5963_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5963_2_i) );
// C_AND/D//AND/D      x66y61     80'h00_FA00_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5964_1 ( .OUT(na5964_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2590_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5964_2 ( .OUT(na5964_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5964_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5964_4 ( .OUT(na5964_2_i), .IN1(na2562_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5964_5 ( .OUT(na5964_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5964_2_i) );
// C_AND/D//AND/D      x66y55     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5965_1 ( .OUT(na5965_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2592_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5965_2 ( .OUT(na5965_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5965_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5965_4 ( .OUT(na5965_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2563_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5965_5 ( .OUT(na5965_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5965_2_i) );
// C_AND/D//AND/D      x63y69     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5967_1 ( .OUT(na5967_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2568_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5967_2 ( .OUT(na5967_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5967_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5967_4 ( .OUT(na5967_2_i), .IN1(1'b1), .IN2(na2567_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5967_5 ( .OUT(na5967_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5967_2_i) );
// C_AND/D//AND/D      x66y76     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5969_1 ( .OUT(na5969_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2570_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5969_2 ( .OUT(na5969_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5969_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5969_4 ( .OUT(na5969_2_i), .IN1(na2569_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5969_5 ( .OUT(na5969_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5969_2_i) );
// C_AND/D//AND/D      x63y77     80'h00_FA00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5971_1 ( .OUT(na5971_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2572_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5971_2 ( .OUT(na5971_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5971_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5971_4 ( .OUT(na5971_2_i), .IN1(1'b1), .IN2(na2571_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5971_5 ( .OUT(na5971_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5971_2_i) );
// C_AND/D///      x51y49     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5972_1 ( .OUT(na5972_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2573_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5972_2 ( .OUT(na5972_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5972_1_i) );
// C_///AND/D      x78y58     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5974_4 ( .OUT(na5974_2_i), .IN1(1'b1), .IN2(na5977_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5974_5 ( .OUT(na5974_2), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5974_2_i) );
// C_AND/D///      x73y76     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5977_1 ( .OUT(na5977_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3325_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5977_2 ( .OUT(na5977_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5977_1_i) );
// C_AND/D///      x63y50     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5985_1 ( .OUT(na5985_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1383_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5985_2 ( .OUT(na5985_1), .CLK(na4116_1), .EN(~na406_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na5985_1_i) );
// C_AND/D///      x87y113     80'h00_D900_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6004_1 ( .OUT(na6004_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2732_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6004_2 ( .OUT(na6004_1), .CLK(~na4116_1), .EN(na3593_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6004_1_i) );
// C_///AND/D      x102y96     80'h00_D900_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6005_4 ( .OUT(na6005_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6047_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6005_5 ( .OUT(na6005_2), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6005_2_i) );
// C_AND/D///      x120y112     80'h00_D900_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6006_1 ( .OUT(na6006_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6047_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6006_2 ( .OUT(na6006_1), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6006_1_i) );
// C_///AND/D      x126y108     80'h00_D900_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6007_4 ( .OUT(na6007_2_i), .IN1(1'b1), .IN2(na6049_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6007_5 ( .OUT(na6007_2), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6007_2_i) );
// C_AND/D///      x122y115     80'h00_D900_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6008_1 ( .OUT(na6008_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6049_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6008_2 ( .OUT(na6008_1), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6008_1_i) );
// C_///AND/D      x122y115     80'h00_D900_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6009_4 ( .OUT(na6009_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6051_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6009_5 ( .OUT(na6009_2), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6009_2_i) );
// C_AND/D///      x123y120     80'h00_D900_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6010_1 ( .OUT(na6010_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6051_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6010_2 ( .OUT(na6010_1), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6010_1_i) );
// C_///AND/D      x122y113     80'h00_D900_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6011_4 ( .OUT(na6011_2_i), .IN1(1'b1), .IN2(na6053_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6011_5 ( .OUT(na6011_2), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6011_2_i) );
// C_AND/D///      x121y115     80'h00_D900_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6012_1 ( .OUT(na6012_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6053_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6012_2 ( .OUT(na6012_1), .CLK(~na4116_1), .EN(na3240_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6012_1_i) );
// C_///AND/D      x86y70     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6014_4 ( .OUT(na6014_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1904_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6014_5 ( .OUT(na6014_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6014_2_i) );
// C_AND/D///      x86y70     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6015_1 ( .OUT(na6015_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1922_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6015_2 ( .OUT(na6015_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6015_1_i) );
// C_///AND/D      x84y82     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6016_4 ( .OUT(na6016_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1932_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6016_5 ( .OUT(na6016_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6016_2_i) );
// C_AND/D///      x80y79     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6017_1 ( .OUT(na6017_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1942_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6017_2 ( .OUT(na6017_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6017_1_i) );
// C_///AND/D      x83y71     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6018_4 ( .OUT(na6018_2_i), .IN1(1'b1), .IN2(na1951_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6018_5 ( .OUT(na6018_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6018_2_i) );
// C_AND/D///      x89y56     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6019_1 ( .OUT(na6019_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1960_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6019_2 ( .OUT(na6019_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6019_1_i) );
// C_///AND/D      x79y77     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6020_4 ( .OUT(na6020_2_i), .IN1(1'b1), .IN2(na1969_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6020_5 ( .OUT(na6020_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6020_2_i) );
// C_AND/D///      x87y72     80'h00_F600_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6021_1 ( .OUT(na6021_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1978_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6021_2 ( .OUT(na6021_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6021_1_i) );
// C_///AND/D      x102y43     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6022_4 ( .OUT(na6022_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1987_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6022_5 ( .OUT(na6022_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6022_2_i) );
// C_AND/D///      x78y61     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6023_1 ( .OUT(na6023_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1994_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6023_2 ( .OUT(na6023_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6023_1_i) );
// C_///AND/D      x100y41     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6024_4 ( .OUT(na6024_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2001_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6024_5 ( .OUT(na6024_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6024_2_i) );
// C_AND/D///      x83y51     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6025_1 ( .OUT(na6025_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2008_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6025_2 ( .OUT(na6025_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6025_1_i) );
// C_///AND/D      x86y49     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6026_4 ( .OUT(na6026_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2015_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6026_5 ( .OUT(na6026_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6026_2_i) );
// C_AND/D///      x87y58     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6027_1 ( .OUT(na6027_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2022_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6027_2 ( .OUT(na6027_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6027_1_i) );
// C_///AND/D      x86y53     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6028_4 ( .OUT(na6028_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2029_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6028_5 ( .OUT(na6028_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6028_2_i) );
// C_AND/D///      x83y63     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6029_1 ( .OUT(na6029_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2036_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6029_2 ( .OUT(na6029_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6029_1_i) );
// C_///AND/D      x85y71     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6030_4 ( .OUT(na6030_2_i), .IN1(1'b1), .IN2(na2043_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6030_5 ( .OUT(na6030_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6030_2_i) );
// C_AND/D///      x85y51     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6031_1 ( .OUT(na6031_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2050_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6031_2 ( .OUT(na6031_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6031_1_i) );
// C_///AND/D      x83y69     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6032_4 ( .OUT(na6032_2_i), .IN1(1'b1), .IN2(na2057_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6032_5 ( .OUT(na6032_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6032_2_i) );
// C_AND/D///      x86y53     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6033_1 ( .OUT(na6033_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2064_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6033_2 ( .OUT(na6033_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6033_1_i) );
// C_///AND/D      x87y69     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6034_4 ( .OUT(na6034_2_i), .IN1(1'b1), .IN2(na2071_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6034_5 ( .OUT(na6034_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6034_2_i) );
// C_AND/D///      x86y55     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6035_1 ( .OUT(na6035_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2078_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6035_2 ( .OUT(na6035_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6035_1_i) );
// C_///AND/D      x83y63     80'h00_F600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6036_4 ( .OUT(na6036_2_i), .IN1(1'b1), .IN2(na2085_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6036_5 ( .OUT(na6036_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6036_2_i) );
// C_AND/D///      x87y53     80'h00_F600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6037_1 ( .OUT(na6037_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2092_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6037_2 ( .OUT(na6037_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6037_1_i) );
// C_///AND/D      x112y45     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6038_4 ( .OUT(na6038_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2099_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6038_5 ( .OUT(na6038_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6038_2_i) );
// C_AND/D///      x88y57     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6039_1 ( .OUT(na6039_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2106_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6039_2 ( .OUT(na6039_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6039_1_i) );
// C_///AND/D      x90y55     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6040_4 ( .OUT(na6040_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2113_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6040_5 ( .OUT(na6040_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6040_2_i) );
// C_AND/D///      x90y59     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6041_1 ( .OUT(na6041_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2120_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6041_2 ( .OUT(na6041_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6041_1_i) );
// C_///AND/D      x100y53     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6042_4 ( .OUT(na6042_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2127_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6042_5 ( .OUT(na6042_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6042_2_i) );
// C_AND/D///      x90y57     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6043_1 ( .OUT(na6043_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2134_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6043_2 ( .OUT(na6043_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6043_1_i) );
// C_///AND/D      x88y55     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6044_4 ( .OUT(na6044_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2141_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6044_5 ( .OUT(na6044_2), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6044_2_i) );
// C_AND/D///      x86y61     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6045_1 ( .OUT(na6045_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2148_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6045_2 ( .OUT(na6045_1), .CLK(na4116_1), .EN(~na340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6045_1_i) );
// C_AND/D//AND/D      x122y123     80'h00_F900_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6047_1 ( .OUT(na6047_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6611_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6047_2 ( .OUT(na6047_1), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6047_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6047_4 ( .OUT(na6047_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6047_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6047_5 ( .OUT(na6047_2), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6047_2_i) );
// C_AND/D//AND/D      x123y122     80'h00_F900_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6049_1 ( .OUT(na6049_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6047_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6049_2 ( .OUT(na6049_1), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6049_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6049_4 ( .OUT(na6049_2_i), .IN1(1'b1), .IN2(na6049_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6049_5 ( .OUT(na6049_2), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6049_2_i) );
// C_AND/D//AND/D      x122y122     80'h00_F900_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6051_1 ( .OUT(na6051_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6049_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6051_2 ( .OUT(na6051_1), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6051_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6051_4 ( .OUT(na6051_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6051_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6051_5 ( .OUT(na6051_2), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6051_2_i) );
// C_AND/D//AND/D      x121y122     80'h00_F900_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6053_1 ( .OUT(na6053_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6051_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6053_2 ( .OUT(na6053_1), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6053_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6053_4 ( .OUT(na6053_2_i), .IN1(1'b1), .IN2(na6053_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6053_5 ( .OUT(na6053_2), .CLK(~na4116_1), .EN(na3234_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6053_2_i) );
// C_AND/D//AND/D      x127y113     80'h00_F900_80_0000_0C88_F5FA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6055_1 ( .OUT(na6055_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2693_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6055_2 ( .OUT(na6055_1), .CLK(~na4116_1), .EN(na3232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6055_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6055_4 ( .OUT(na6055_2_i), .IN1(na2693_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6055_5 ( .OUT(na6055_2), .CLK(~na4116_1), .EN(na3232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6055_2_i) );
// C_/C_0_1///      x83y103     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a6056_2 ( .OUT(na6056_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a6056_6 ( .COUTY1(na6056_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6056_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND/L///      x104y115     80'h10_DE00_00_0000_0C88_FFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6057_1 ( .OUT(na6057_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_L        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6057_2 ( .OUT(na6057_1), .CLK(na3_1), .EN(1'b1), .SR(~na1_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6057_1_i) );
// C_///AND/L      x76y35     80'h10_DE00_80_0000_0C08_FFFF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6058_4 ( .OUT(na6058_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_L        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6058_5 ( .OUT(na6058_2), .CLK(na4_2), .EN(1'b1), .SR(~na2_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6058_2_i) );
// C_///AND/D      x117y102     80'h00_DD00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6065_4 ( .OUT(na6065_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2734_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6065_5 ( .OUT(na6065_2), .CLK(~na4116_1), .EN(1'b1), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6065_2_i) );
// C_AND/D///      x130y99     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6066_1 ( .OUT(na6066_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3214_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6066_2 ( .OUT(na6066_1), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6066_1_i) );
// C_///AND/D      x104y101     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6067_4 ( .OUT(na6067_2_i), .IN1(na3494_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6067_5 ( .OUT(na6067_2), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6067_2_i) );
// C_AND/D///      x125y110     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6068_1 ( .OUT(na6068_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na107_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6068_2 ( .OUT(na6068_1), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6068_1_i) );
// C_///AND/D      x125y102     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6069_4 ( .OUT(na6069_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na116_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6069_5 ( .OUT(na6069_2), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6069_2_i) );
// C_AND/D///      x122y109     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6070_1 ( .OUT(na6070_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3496_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6070_2 ( .OUT(na6070_1), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6070_1_i) );
// C_///AND/D      x124y111     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6071_4 ( .OUT(na6071_2_i), .IN1(na129_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6071_5 ( .OUT(na6071_2), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6071_2_i) );
// C_AND/D///      x125y115     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6072_1 ( .OUT(na6072_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na135_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6072_2 ( .OUT(na6072_1), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6072_1_i) );
// C_///AND/D      x126y110     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6073_4 ( .OUT(na6073_2_i), .IN1(1'b1), .IN2(na142_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6073_5 ( .OUT(na6073_2), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6073_2_i) );
// C_AND/D///      x125y119     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6074_1 ( .OUT(na6074_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na149_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6074_2 ( .OUT(na6074_1), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6074_1_i) );
// C_///AND/D      x118y99     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6075_4 ( .OUT(na6075_2_i), .IN1(na3258_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6075_5 ( .OUT(na6075_2), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6075_2_i) );
// C_AND/D///      x119y102     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6076_1 ( .OUT(na6076_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3499_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6076_2 ( .OUT(na6076_1), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6076_1_i) );
// C_///AND/D      x128y115     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6077_4 ( .OUT(na6077_2_i), .IN1(na103_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6077_5 ( .OUT(na6077_2), .CLK(na4116_1), .EN(na3340_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6077_2_i) );
// C_AND/D///      x128y102     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6078_1 ( .OUT(na6078_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3214_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6078_2 ( .OUT(na6078_1), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6078_1_i) );
// C_///AND/D      x128y120     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6079_4 ( .OUT(na6079_2_i), .IN1(na3494_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6079_5 ( .OUT(na6079_2), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6079_2_i) );
// C_AND/D///      x123y111     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6080_1 ( .OUT(na6080_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na107_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6080_2 ( .OUT(na6080_1), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6080_1_i) );
// C_///AND/D      x125y107     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6081_4 ( .OUT(na6081_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na116_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6081_5 ( .OUT(na6081_2), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6081_2_i) );
// C_AND/D///      x122y112     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6082_1 ( .OUT(na6082_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3496_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6082_2 ( .OUT(na6082_1), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6082_1_i) );
// C_///AND/D      x124y112     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6083_4 ( .OUT(na6083_2_i), .IN1(na129_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6083_5 ( .OUT(na6083_2), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6083_2_i) );
// C_AND/D///      x125y116     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6084_1 ( .OUT(na6084_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na135_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6084_2 ( .OUT(na6084_1), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6084_1_i) );
// C_///AND/D      x126y111     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6085_4 ( .OUT(na6085_2_i), .IN1(1'b1), .IN2(na142_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6085_5 ( .OUT(na6085_2), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6085_2_i) );
// C_AND/D///      x127y120     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6086_1 ( .OUT(na6086_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na149_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6086_2 ( .OUT(na6086_1), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6086_1_i) );
// C_///AND/D      x118y98     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6087_4 ( .OUT(na6087_2_i), .IN1(na3258_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6087_5 ( .OUT(na6087_2), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6087_2_i) );
// C_AND/D///      x115y99     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6088_1 ( .OUT(na6088_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3499_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6088_2 ( .OUT(na6088_1), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6088_1_i) );
// C_///AND/D      x136y116     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6089_4 ( .OUT(na6089_2_i), .IN1(na103_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6089_5 ( .OUT(na6089_2), .CLK(na4116_1), .EN(na3341_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6089_2_i) );
// C_AND/D///      x65y36     80'h00_D500_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6090_1 ( .OUT(na6090_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2758_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6090_2 ( .OUT(na6090_1), .CLK(~na4116_1), .EN(~na3253_1), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6090_1_i) );
// C_///AND/D      x125y56     80'h00_D900_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6091_4 ( .OUT(na6091_2_i), .IN1(1'b1), .IN2(na6105_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6091_5 ( .OUT(na6091_2), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6091_2_i) );
// C_AND/D///      x120y64     80'h00_D900_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6092_1 ( .OUT(na6092_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6105_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6092_2 ( .OUT(na6092_1), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6092_1_i) );
// C_///AND/D      x130y56     80'h00_D900_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6093_4 ( .OUT(na6093_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6107_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6093_5 ( .OUT(na6093_2), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6093_2_i) );
// C_AND/D///      x127y63     80'h00_D900_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6094_1 ( .OUT(na6094_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6107_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6094_2 ( .OUT(na6094_1), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6094_1_i) );
// C_///AND/D      x132y60     80'h00_D900_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6095_4 ( .OUT(na6095_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6109_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6095_5 ( .OUT(na6095_2), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6095_2_i) );
// C_AND/D///      x132y68     80'h00_D900_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6096_1 ( .OUT(na6096_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6109_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6096_2 ( .OUT(na6096_1), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6096_1_i) );
// C_///AND/D      x129y62     80'h00_D900_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6097_4 ( .OUT(na6097_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6111_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6097_5 ( .OUT(na6097_2), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6097_2_i) );
// C_AND/D///      x132y70     80'h00_D900_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6098_1 ( .OUT(na6098_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6111_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6098_2 ( .OUT(na6098_1), .CLK(~na4116_1), .EN(na3274_2), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6098_1_i) );
// C_AND/D//AND/D      x129y64     80'h00_F900_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6105_1 ( .OUT(na6105_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6607_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6105_2 ( .OUT(na6105_1), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6105_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6105_4 ( .OUT(na6105_2_i), .IN1(1'b1), .IN2(na6105_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6105_5 ( .OUT(na6105_2), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6105_2_i) );
// C_AND/D//AND/D      x130y63     80'h00_F900_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6107_1 ( .OUT(na6107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6105_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6107_2 ( .OUT(na6107_1), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6107_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6107_4 ( .OUT(na6107_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6107_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6107_5 ( .OUT(na6107_2), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6107_2_i) );
// C_AND/D//AND/D      x134y64     80'h00_F900_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6109_1 ( .OUT(na6109_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na6107_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6109_2 ( .OUT(na6109_1), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6109_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6109_4 ( .OUT(na6109_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na6109_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6109_5 ( .OUT(na6109_2), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6109_2_i) );
// C_AND/D//AND/D      x132y63     80'h00_F900_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6111_1 ( .OUT(na6111_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6109_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6111_2 ( .OUT(na6111_1), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6111_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6111_4 ( .OUT(na6111_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na6111_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a6111_5 ( .OUT(na6111_2), .CLK(~na4116_1), .EN(na3251_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6111_2_i) );
// C_///AND/D      x121y44     80'h00_F900_80_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6113_4 ( .OUT(na6113_2_i), .IN1(~na2832_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6113_5 ( .OUT(na6113_2), .CLK(~na4116_1), .EN(na3250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6113_2_i) );
// C_AND/D///      x118y50     80'h00_F900_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6117_1 ( .OUT(na6117_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2832_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6117_2 ( .OUT(na6117_1), .CLK(~na4116_1), .EN(na3250_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6117_1_i) );
// C_///AND/D      x105y65     80'h00_DD00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6118_4 ( .OUT(na6118_2_i), .IN1(1'b1), .IN2(na2760_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6118_5 ( .OUT(na6118_2), .CLK(~na4116_1), .EN(1'b1), .SR(~na6626_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6118_2_i) );
// C_AND/D///      x60y79     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6308_1 ( .OUT(na6308_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5795_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6308_2 ( .OUT(na6308_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6308_1_i) );
// C_///AND/D      x72y86     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6309_4 ( .OUT(na6309_2_i), .IN1(1'b1), .IN2(na5796_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6309_5 ( .OUT(na6309_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6309_2_i) );
// C_AND/D///      x56y80     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6310_1 ( .OUT(na6310_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5797_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6310_2 ( .OUT(na6310_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6310_1_i) );
// C_///AND/D      x51y79     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6312_4 ( .OUT(na6312_2_i), .IN1(na5799_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6312_5 ( .OUT(na6312_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6312_2_i) );
// C_AND/D///      x51y79     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6313_1 ( .OUT(na6313_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5800_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6313_2 ( .OUT(na6313_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6313_1_i) );
// C_///AND/D      x50y79     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6314_4 ( .OUT(na6314_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5801_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6314_5 ( .OUT(na6314_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6314_2_i) );
// C_AND/D///      x51y77     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6315_1 ( .OUT(na6315_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5802_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6315_2 ( .OUT(na6315_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6315_1_i) );
// C_///AND/D      x53y77     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6317_4 ( .OUT(na6317_2_i), .IN1(na5804_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6317_5 ( .OUT(na6317_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6317_2_i) );
// C_AND/D///      x49y79     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6318_1 ( .OUT(na6318_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5805_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6318_2 ( .OUT(na6318_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6318_1_i) );
// C_///AND/D      x49y75     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6319_4 ( .OUT(na6319_2_i), .IN1(na5806_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6319_5 ( .OUT(na6319_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6319_2_i) );
// C_AND/D//AND/D      x49y83     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6320_1 ( .OUT(na6320_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5807_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6320_2 ( .OUT(na6320_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6320_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6320_4 ( .OUT(na6320_2_i), .IN1(1'b1), .IN2(na5824_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6320_5 ( .OUT(na6320_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6320_2_i) );
// C_AND/D///      x51y75     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6321_1 ( .OUT(na6321_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5808_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6321_2 ( .OUT(na6321_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6321_1_i) );
// C_///AND/D      x51y75     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6322_4 ( .OUT(na6322_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5809_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6322_5 ( .OUT(na6322_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6322_2_i) );
// C_AND/D///      x53y77     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6323_1 ( .OUT(na6323_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5810_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6323_2 ( .OUT(na6323_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6323_1_i) );
// C_AND/D//AND/D      x53y75     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6324_1 ( .OUT(na6324_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5811_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6324_2 ( .OUT(na6324_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6324_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6324_4 ( .OUT(na6324_2_i), .IN1(1'b1), .IN2(na5798_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6324_5 ( .OUT(na6324_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6324_2_i) );
// C_AND/D//AND/D      x49y77     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6325_1 ( .OUT(na6325_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5812_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6325_2 ( .OUT(na6325_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6325_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6325_4 ( .OUT(na6325_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5803_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6325_5 ( .OUT(na6325_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6325_2_i) );
// C_///AND/D      x65y93     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6326_4 ( .OUT(na6326_2_i), .IN1(1'b1), .IN2(na5813_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6326_5 ( .OUT(na6326_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6326_2_i) );
// C_AND/D///      x55y77     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6327_1 ( .OUT(na6327_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5814_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6327_2 ( .OUT(na6327_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6327_1_i) );
// C_///AND/D      x67y89     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6328_4 ( .OUT(na6328_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5815_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6328_5 ( .OUT(na6328_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6328_2_i) );
// C_AND/D///      x58y79     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6329_1 ( .OUT(na6329_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5816_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6329_2 ( .OUT(na6329_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6329_1_i) );
// C_///AND/D      x58y79     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6330_4 ( .OUT(na6330_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5817_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6330_5 ( .OUT(na6330_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6330_2_i) );
// C_AND/D///      x51y81     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6331_1 ( .OUT(na6331_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5818_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6331_2 ( .OUT(na6331_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6331_1_i) );
// C_///AND/D      x67y91     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6332_4 ( .OUT(na6332_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5819_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6332_5 ( .OUT(na6332_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6332_2_i) );
// C_AND/D///      x47y81     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6333_1 ( .OUT(na6333_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na5820_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6333_2 ( .OUT(na6333_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6333_1_i) );
// C_///AND/D      x51y77     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6334_4 ( .OUT(na6334_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5821_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6334_5 ( .OUT(na6334_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6334_2_i) );
// C_AND/D///      x49y81     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6335_1 ( .OUT(na6335_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na5822_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6335_2 ( .OUT(na6335_1), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6335_1_i) );
// C_///AND/D      x67y81     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6336_4 ( .OUT(na6336_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5823_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6336_5 ( .OUT(na6336_2), .CLK(na4116_1), .EN(na504_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6336_2_i) );
// C_ADDF////      x54y60     80'h00_0018_00_0010_0666_00AC
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a6343_1 ( .OUT(na6343_1), .COUTY1(na6343_4), .IN1(1'b1), .IN2(na3598_2), .IN3(na357_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na2627_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y66     80'h00_0078_00_0020_0C66_A9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6345_1 ( .OUT(na6345_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2378_2), .IN6(na3598_2), .IN7(na2316_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6374_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6345_4 ( .OUT(na6345_2), .COUTY1(na6345_4), .IN1(~na2378_1), .IN2(na3598_2), .IN3(na607_1), .IN4(1'b0), .IN5(~na2378_2),
                      .IN6(na3598_2), .IN7(na2316_2), .IN8(1'b0), .CINX(1'b0), .CINY1(na6374_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y67     80'h00_0078_00_0020_0C66_C9C9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6347_1 ( .OUT(na6347_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9586_2), .IN6(na3598_2), .IN7(1'b0), .IN8(na612_1),
                      .CINX(1'b0), .CINY1(na6345_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6347_4 ( .OUT(na6347_2), .COUTY1(na6347_4), .IN1(~na2354_1), .IN2(na3598_2), .IN3(1'b0), .IN4(na622_1), .IN5(~na9586_2),
                      .IN6(na3598_2), .IN7(1'b0), .IN8(na612_1), .CINX(1'b0), .CINY1(na6345_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y68     80'h00_0078_00_0020_0C66_C9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6349_1 ( .OUT(na6349_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2383_2), .IN6(na3598_2), .IN7(1'b0), .IN8(na617_1),
                      .CINX(1'b0), .CINY1(na6347_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6349_4 ( .OUT(na6349_2), .COUTY1(na6349_4), .IN1(~na2383_1), .IN2(na3598_2), .IN3(na627_1), .IN4(1'b0), .IN5(~na2383_2),
                      .IN6(na3598_2), .IN7(1'b0), .IN8(na617_1), .CINX(1'b0), .CINY1(na6347_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y69     80'h00_0078_00_0020_0C66_A9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6351_1 ( .OUT(na6351_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9587_2), .IN6(na3598_2), .IN7(na9526_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6349_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6351_4 ( .OUT(na6351_2), .COUTY1(na6351_4), .IN1(~na9590_2), .IN2(na3598_2), .IN3(na632_1), .IN4(1'b0), .IN5(~na9587_2),
                      .IN6(na3598_2), .IN7(na9526_2), .IN8(1'b0), .CINX(1'b0), .CINY1(na6349_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y70     80'h00_0078_00_0020_0C66_A9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6353_1 ( .OUT(na6353_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2332_1), .IN6(na3598_2), .IN7(na637_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6351_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6353_4 ( .OUT(na6353_2), .COUTY1(na6353_4), .IN1(~na9585_2), .IN2(na3598_2), .IN3(na9522_2), .IN4(1'b0), .IN5(~na2332_1),
                      .IN6(na3598_2), .IN7(na637_1), .IN8(1'b0), .CINX(1'b0), .CINY1(na6351_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y61     80'h00_0078_00_0020_0C66_C9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6354_1 ( .OUT(na6354_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na50_2), .IN6(na3598_2), .IN7(1'b0), .IN8(na355_1),
                      .CINX(1'b0), .CINY1(na6343_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6354_4 ( .OUT(na6354_2), .COUTY1(na6354_4), .IN1(~na9825_2), .IN2(na3598_2), .IN3(na9253_2), .IN4(1'b0), .IN5(~na50_2), .IN6(na3598_2),
                      .IN7(1'b0), .IN8(na355_1), .CINX(1'b0), .CINY1(na6343_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y71     80'h00_0078_00_0020_0C66_A9C9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6356_1 ( .OUT(na6356_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9570_2), .IN6(na3598_2), .IN7(na661_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6353_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6356_4 ( .OUT(na6356_2), .COUTY1(na6356_4), .IN1(~na9571_2), .IN2(na3598_2), .IN3(1'b0), .IN4(na667_1), .IN5(~na9570_2),
                      .IN6(na3598_2), .IN7(na661_1), .IN8(1'b0), .CINX(1'b0), .CINY1(na6353_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y72     80'h00_0078_00_0020_0C66_A9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6358_1 ( .OUT(na6358_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2351_2), .IN6(na3598_2), .IN7(na672_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6356_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6358_4 ( .OUT(na6358_2), .COUTY1(na6358_4), .IN1(~na9584_2), .IN2(na3598_2), .IN3(na677_1), .IN4(1'b0), .IN5(~na2351_2),
                      .IN6(na3598_2), .IN7(na672_1), .IN8(1'b0), .CINX(1'b0), .CINY1(na6356_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y73     80'h00_0078_00_0020_0C66_C9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6360_1 ( .OUT(na6360_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9582_2), .IN6(na3598_2), .IN7(1'b0), .IN8(na682_1),
                      .CINX(1'b0), .CINY1(na6358_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6360_4 ( .OUT(na6360_2), .COUTY1(na6360_4), .IN1(~na9575_2), .IN2(na3598_2), .IN3(na9310_2), .IN4(1'b0), .IN5(~na9582_2),
                      .IN6(na3598_2), .IN7(1'b0), .IN8(na682_1), .CINX(1'b0), .CINY1(na6358_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y74     80'h00_0078_00_0020_0C66_A9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6362_1 ( .OUT(na6362_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9569_2), .IN6(na3598_2), .IN7(na692_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6360_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6362_4 ( .OUT(na6362_2), .COUTY1(na6362_4), .IN1(~na2309_1), .IN2(na3598_2), .IN3(na9315_2), .IN4(1'b0), .IN5(~na9569_2),
                      .IN6(na3598_2), .IN7(na692_1), .IN8(1'b0), .CINX(1'b0), .CINY1(na6360_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y75     80'h00_0078_00_0020_0C66_C9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6364_1 ( .OUT(na6364_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2385_1), .IN6(na3598_2), .IN7(1'b0), .IN8(na702_1),
                      .CINX(1'b0), .CINY1(na6362_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6364_4 ( .OUT(na6364_2), .COUTY1(na6364_4), .IN1(~na2351_1), .IN2(na3598_2), .IN3(na707_1), .IN4(1'b0), .IN5(~na2385_1),
                      .IN6(na3598_2), .IN7(1'b0), .IN8(na702_1), .CINX(1'b0), .CINY1(na6362_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDFx////      x54y76     80'h00_0018_00_0010_0666_00A9
C_ADDFx    #(.CPE_CFG (9'b0_0010_0000)) 
           _a6367_1 ( .OUT(na6367_1), .IN1(~na2354_2), .IN2(na3598_2), .IN3(na723_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6364_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y62     80'h00_0078_00_0020_0C66_A9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6368_1 ( .OUT(na6368_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9824_2), .IN6(na3598_2), .IN7(na545_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6354_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6368_4 ( .OUT(na6368_2), .COUTY1(na6368_4), .IN1(~na3487_1), .IN2(na3598_2), .IN3(na550_1), .IN4(1'b0), .IN5(~na9824_2),
                      .IN6(na3598_2), .IN7(na545_1), .IN8(1'b0), .CINX(1'b0), .CINY1(na6354_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y63     80'h00_0078_00_0020_0C66_A9C9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6370_1 ( .OUT(na6370_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9592_2), .IN6(na3598_2), .IN7(na2369_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6368_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6370_4 ( .OUT(na6370_2), .COUTY1(na6370_4), .IN1(~na2362_1), .IN2(na3598_2), .IN3(1'b0), .IN4(na2348_2), .IN5(~na9592_2),
                      .IN6(na3598_2), .IN7(na2369_2), .IN8(1'b0), .CINX(1'b0), .CINY1(na6368_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y64     80'h00_0078_00_0020_0C66_A9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6372_1 ( .OUT(na6372_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9275_2), .IN6(na3598_2), .IN7(na9568_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(na6370_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6372_4 ( .OUT(na6372_2), .COUTY1(na6372_4), .IN1(~na2338_2), .IN2(na3598_2), .IN3(na589_1), .IN4(1'b0), .IN5(~na9275_2),
                      .IN6(na3598_2), .IN7(na9568_2), .IN8(1'b0), .CINX(1'b0), .CINY1(na6370_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x///ADDF2x/      x54y65     80'h00_0078_00_0020_0C66_C9A9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a6374_1 ( .OUT(na6374_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9580_2), .IN6(na3598_2), .IN7(1'b0), .IN8(na594_1),
                      .CINX(1'b0), .CINY1(na6372_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a6374_4 ( .OUT(na6374_2), .COUTY1(na6374_4), .IN1(~na2332_2), .IN2(na3598_2), .IN3(na2327_2), .IN4(1'b0), .IN5(~na9580_2),
                      .IN6(na3598_2), .IN7(1'b0), .IN8(na594_1), .CINX(1'b0), .CINY1(na6372_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDFx////      x76y124     80'h00_0018_00_0010_0666_00A6
C_ADDFx    #(.CPE_CFG (9'b0_0010_0000)) 
           _a6380_1 ( .OUT(na6380_1), .COUTY1(na6380_4), .IN1(~na3335_2), .IN2(~na713_1), .IN3(na1433_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na6562_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x76y125     80'h00_0078_00_0020_0C66_55A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a6381_1 ( .OUT(na6381_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3421_1), .IN6(1'b1), .IN7(~na1433_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na6380_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a6381_4 ( .OUT(na6381_2), .IN1(1'b1), .IN2(~na1414_2), .IN3(na1433_1), .IN4(1'b1), .IN5(~na3421_1), .IN6(1'b1), .IN7(~na1433_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na6380_4), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y53     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6383_1 ( .OUT(na6383_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9979_2), .IN6(na10003_2), .IN7(na8604_1),
                      .IN8(na10099_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x90y60     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6384_1 ( .OUT(na6384_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10119_2), .IN6(na10163_2), .IN7(na7821_1),
                      .IN8(na10024_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6385_1 ( .OUT(na6385_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9978_2), .IN6(na10002_2), .IN7(na8603_2),
                      .IN8(na10098_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y57     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6386_1 ( .OUT(na6386_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10118_2), .IN6(na10162_2), .IN7(na7819_2),
                      .IN8(na10023_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x71y52     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6387_1 ( .OUT(na6387_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9977_2), .IN6(na10001_2), .IN7(na10073_2),
                      .IN8(na8738_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y51     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6388_1 ( .OUT(na6388_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10117_2), .IN6(na10161_2), .IN7(na9983_2),
                      .IN8(na8038_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x67y52     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6389_1 ( .OUT(na6389_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9976_2), .IN6(na10000_2), .IN7(na10072_2),
                      .IN8(na8737_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y53     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6390_1 ( .OUT(na6390_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10116_2), .IN6(na10160_2), .IN7(na9982_2),
                      .IN8(na8037_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y52     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6391_1 ( .OUT(na6391_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9975_2), .IN6(na9999_2), .IN7(na8600_1),
                      .IN8(na10065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y49     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6392_1 ( .OUT(na6392_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10115_2), .IN6(na10159_2), .IN7(na7809_1),
                      .IN8(na10022_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6393_1 ( .OUT(na6393_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9974_2), .IN6(na9998_2), .IN7(na8599_2),
                      .IN8(na10064_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y51     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6394_1 ( .OUT(na6394_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10114_2), .IN6(na10158_2), .IN7(na7807_2),
                      .IN8(na10021_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y56     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6395_1 ( .OUT(na6395_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9973_2), .IN6(na9997_2), .IN7(na10071_2),
                      .IN8(na8510_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6396_1 ( .OUT(na6396_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10113_2), .IN6(na10157_2), .IN7(na9981_2),
                      .IN8(na8032_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y56     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6397_1 ( .OUT(na6397_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9972_2), .IN6(na9996_2), .IN7(na10070_2),
                      .IN8(na8509_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y53     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6398_1 ( .OUT(na6398_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10112_2), .IN6(na10156_2), .IN7(na9980_2),
                      .IN8(na8031_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y69     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6399_1 ( .OUT(na6399_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9971_2), .IN6(na10097_2), .IN7(na8596_1),
                      .IN8(na10063_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y62     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6400_1 ( .OUT(na6400_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10111_2), .IN6(na10155_2), .IN7(na8199_1),
                      .IN8(na10020_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y73     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6401_1 ( .OUT(na6401_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9970_2), .IN6(na10096_2), .IN7(na8595_2),
                      .IN8(na10062_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x75y66     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6402_1 ( .OUT(na6402_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10110_2), .IN6(na10154_2), .IN7(na8198_2),
                      .IN8(na10019_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y70     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6403_1 ( .OUT(na6403_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9969_2), .IN6(na10095_2), .IN7(na10069_2),
                      .IN8(na8506_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y63     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6404_1 ( .OUT(na6404_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10109_2), .IN6(na10153_2), .IN7(na10039_2),
                      .IN8(na8026_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y72     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6405_1 ( .OUT(na6405_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9968_2), .IN6(na10094_2), .IN7(na10068_2),
                      .IN8(na8505_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y69     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6406_1 ( .OUT(na6406_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10108_2), .IN6(na10152_2), .IN7(na10038_2),
                      .IN8(na8025_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y73     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6407_1 ( .OUT(na6407_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9967_2), .IN6(na10093_2), .IN7(na8592_1),
                      .IN8(na10061_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y56     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6408_1 ( .OUT(na6408_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10143_2), .IN6(na10151_2), .IN7(na8194_1),
                      .IN8(na10018_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y70     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6409_1 ( .OUT(na6409_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9966_2), .IN6(na10092_2), .IN7(na8591_2),
                      .IN8(na10060_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x84y61     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6410_1 ( .OUT(na6410_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10142_2), .IN6(na10150_2), .IN7(na8193_2),
                      .IN8(na10017_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y74     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6411_1 ( .OUT(na6411_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9965_2), .IN6(na10091_2), .IN7(na10067_2),
                      .IN8(na8502_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y61     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6412_1 ( .OUT(na6412_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10141_2), .IN6(na10149_2), .IN7(na10037_2),
                      .IN8(na8020_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y75     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6413_1 ( .OUT(na6413_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9964_2), .IN6(na10090_2), .IN7(na10066_2),
                      .IN8(na8501_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x84y64     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6414_1 ( .OUT(na6414_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10140_2), .IN6(na10148_2), .IN7(na10036_2),
                      .IN8(na8019_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y61     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6415_1 ( .OUT(na6415_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9963_2), .IN6(na10089_2), .IN7(na8756_1),
                      .IN8(na10059_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y60     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6416_1 ( .OUT(na6416_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10139_2), .IN6(na10147_2), .IN7(na8188_1),
                      .IN8(na10048_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y62     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6417_1 ( .OUT(na6417_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9962_2), .IN6(na10088_2), .IN7(na8755_2),
                      .IN8(na10058_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y59     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6418_1 ( .OUT(na6418_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10138_2), .IN6(na10146_2), .IN7(na8181_2),
                      .IN8(na10047_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y61     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6419_1 ( .OUT(na6419_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9961_2), .IN6(na10087_2), .IN7(na10107_2),
                      .IN8(na8498_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y64     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6420_1 ( .OUT(na6420_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10137_2), .IN6(na10145_2), .IN7(na10034_2),
                      .IN8(na8217_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y61     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6421_1 ( .OUT(na6421_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na9960_2), .IN6(na10086_2), .IN7(na10106_2),
                      .IN8(na8497_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x73y64     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6422_1 ( .OUT(na6422_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10136_2), .IN6(na10144_2), .IN7(na10033_2),
                      .IN8(na8216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x62y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6423_1 ( .OUT(na6423_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10015_2), .IN6(na10085_2), .IN7(na8752_1),
                      .IN8(na10056_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x82y57     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6424_1 ( .OUT(na6424_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10135_2), .IN6(na9995_2), .IN7(na8178_1),
                      .IN8(na10046_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y52     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6425_1 ( .OUT(na6425_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10014_2), .IN6(na10084_2), .IN7(na8751_2),
                      .IN8(na10055_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y57     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6426_1 ( .OUT(na6426_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10134_2), .IN6(na9994_2), .IN7(na8172_2),
                      .IN8(na10045_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y53     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6427_1 ( .OUT(na6427_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10013_2), .IN6(na10083_2), .IN7(na10105_2),
                      .IN8(na8376_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x75y60     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6428_1 ( .OUT(na6428_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10133_2), .IN6(na9993_2), .IN7(na10032_2),
                      .IN8(na8213_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y53     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6429_1 ( .OUT(na6429_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10012_2), .IN6(na10082_2), .IN7(na10104_2),
                      .IN8(na8374_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6430_1 ( .OUT(na6430_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10132_2), .IN6(na9992_2), .IN7(na10031_2),
                      .IN8(na8212_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y52     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6431_1 ( .OUT(na6431_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10011_2), .IN6(na10081_2), .IN7(na8748_1),
                      .IN8(na10123_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x75y57     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6432_1 ( .OUT(na6432_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10131_2), .IN6(na9991_2), .IN7(na8169_1),
                      .IN8(na10044_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y53     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6433_1 ( .OUT(na6433_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10010_2), .IN6(na10080_2), .IN7(na8747_2),
                      .IN8(na10122_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x75y58     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6434_1 ( .OUT(na6434_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10130_2), .IN6(na9990_2), .IN7(na8168_2),
                      .IN8(na10043_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6435_1 ( .OUT(na6435_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10009_2), .IN6(na10079_2), .IN7(na10103_2),
                      .IN8(na8838_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y61     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6436_1 ( .OUT(na6436_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10129_2), .IN6(na9989_2), .IN7(na10030_2),
                      .IN8(na8209_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x58y53     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6437_1 ( .OUT(na6437_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10008_2), .IN6(na10078_2), .IN7(na10102_2),
                      .IN8(na8837_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y58     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6438_1 ( .OUT(na6438_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10128_2), .IN6(na9988_2), .IN7(na10029_2),
                      .IN8(na8208_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y56     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6439_1 ( .OUT(na6439_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10007_2), .IN6(na10077_2), .IN7(na8744_1),
                      .IN8(na10121_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y57     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6440_1 ( .OUT(na6440_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10127_2), .IN6(na9987_2), .IN7(na8045_1),
                      .IN8(na10042_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y51     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6441_1 ( .OUT(na6441_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10006_2), .IN6(na10076_2), .IN7(na8743_2),
                      .IN8(na10120_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x84y56     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6442_1 ( .OUT(na6442_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10126_2), .IN6(na9986_2), .IN7(na8044_2),
                      .IN8(na10041_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y44     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6443_1 ( .OUT(na6443_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10005_2), .IN6(na10075_2), .IN7(na10101_2),
                      .IN8(na8834_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y59     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6444_1 ( .OUT(na6444_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10125_2), .IN6(na9985_2), .IN7(na10026_2),
                      .IN8(na8205_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y42     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6445_1 ( .OUT(na6445_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10004_2), .IN6(na10074_2), .IN7(na10100_2),
                      .IN8(na8833_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y57     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6446_1 ( .OUT(na6446_1), .IN1(na88_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9163_2), .IN5(na10124_2), .IN6(na9984_2), .IN7(na10025_2),
                      .IN8(na8204_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x98y52     80'h00_FA00_00_0040_0C05_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6447_1 ( .OUT(na6447_1_i), .IN1(na6448_1), .IN2(1'b0), .IN3(na9132_1), .IN4(1'b0), .IN5(1'b1), .IN6(~na59_1), .IN7(1'b1),
                      .IN8(~na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6447_2 ( .OUT(na6447_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6447_1_i) );
// C_MX4a/D///      x93y49     80'h00_FA00_00_0040_0C05_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6448_1 ( .OUT(na6448_1_i), .IN1(na6449_1), .IN2(1'b0), .IN3(na9131_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na59_1), .IN7(1'b1),
                      .IN8(~na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6448_2 ( .OUT(na6448_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6448_1_i) );
// C_MX4a/D///      x93y51     80'h00_FA00_00_0040_0C0A_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6449_1 ( .OUT(na6449_1_i), .IN1(1'b0), .IN2(na6450_1), .IN3(1'b0), .IN4(na9130_1), .IN5(1'b1), .IN6(na59_1), .IN7(1'b1),
                      .IN8(~na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6449_2 ( .OUT(na6449_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6449_1_i) );
// C_MX4a/D///      x93y50     80'h00_FA00_00_0040_0C0A_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6450_1 ( .OUT(na6450_1_i), .IN1(1'b0), .IN2(na6451_1), .IN3(1'b0), .IN4(na9129_2), .IN5(1'b1), .IN6(na59_1), .IN7(1'b1),
                      .IN8(~na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6450_2 ( .OUT(na6450_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6450_1_i) );
// C_MX4a/D///      x93y52     80'h00_FA00_00_0040_0C05_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6451_1 ( .OUT(na6451_1_i), .IN1(na6452_1), .IN2(1'b0), .IN3(na9128_1), .IN4(1'b0), .IN5(1'b1), .IN6(~na59_1), .IN7(1'b1),
                      .IN8(~na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6451_2 ( .OUT(na6451_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6451_1_i) );
// C_MX4a/D///      x93y53     80'h00_FA00_00_0040_0C05_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6452_1 ( .OUT(na6452_1_i), .IN1(na6453_1), .IN2(1'b0), .IN3(na9127_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na59_1), .IN7(1'b1),
                      .IN8(~na973_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6452_2 ( .OUT(na6452_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6452_1_i) );
// C_MX4a/D///      x97y51     80'h00_FA00_00_0040_0C0A_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6453_1 ( .OUT(na6453_1_i), .IN1(1'b0), .IN2(na58_1), .IN3(1'b0), .IN4(na9126_1), .IN5(1'b1), .IN6(na59_1), .IN7(1'b1), .IN8(~na973_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a6453_2 ( .OUT(na6453_1), .CLK(na4116_1), .EN(na59_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6453_1_i) );
// C_MX4b////      x103y61     80'h00_0018_00_0040_0AFC_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6454_1 ( .OUT(na6454_1), .IN1(~na9947_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9146_2), .IN5(na9147_2), .IN6(na9945_2), .IN7(~na76_2),
                      .IN8(~na6673_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x102y67     80'h00_FE00_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6455_1 ( .OUT(na6455_1_i), .IN1(1'b1), .IN2(na67_2), .IN3(na478_2), .IN4(1'b1), .IN5(na6454_1), .IN6(na64_1), .IN7(na478_1),
                      .IN8(na9155_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6455_2 ( .OUT(na6455_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6455_1_i) );
// C_MX4a////      x103y67     80'h00_0018_00_0040_0C4E_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6456_1 ( .OUT(na6456_1), .IN1(1'b0), .IN2(na36_2), .IN3(~na9158_2), .IN4(na73_1), .IN5(na9947_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na9146_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x110y43     80'h00_FE00_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6457_1 ( .OUT(na6457_1_i), .IN1(1'b1), .IN2(na67_2), .IN3(na478_2), .IN4(1'b1), .IN5(na6456_1), .IN6(na69_1), .IN7(na71_1),
                      .IN8(na70_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6457_2 ( .OUT(na6457_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6457_1_i) );
// C_MX4b/D///      x106y63     80'h00_FE00_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6458_1 ( .OUT(na6458_1_i), .IN1(1'b1), .IN2(na67_2), .IN3(na478_2), .IN4(1'b1), .IN5(na72_1), .IN6(na74_1), .IN7(na478_1),
                      .IN8(na75_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6458_2 ( .OUT(na6458_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6458_1_i) );
// C_MX4b////      x102y65     80'h00_0018_00_0040_0AE8_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6459_1 ( .OUT(na6459_1), .IN1(~na9947_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na9146_2), .IN5(1'b0), .IN6(na36_2), .IN7(na76_2),
                      .IN8(~na9149_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y66     80'h00_0018_00_0040_0A90_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6460_1 ( .OUT(na6460_1), .IN1(~na9947_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na9146_2), .IN5(na68_2), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na73_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x114y47     80'h00_FE00_00_0040_0AF0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6461_1 ( .OUT(na6461_1_i), .IN1(1'b1), .IN2(na67_2), .IN3(~na478_2), .IN4(1'b1), .IN5(na77_2), .IN6(na78_1), .IN7(na6459_1),
                      .IN8(na6460_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6461_2 ( .OUT(na6461_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6461_1_i) );
// C_MX4b/D///      x114y46     80'h00_FE00_00_0040_0AF3_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6462_1 ( .OUT(na6462_1_i), .IN1(1'b1), .IN2(na67_2), .IN3(~na478_2), .IN4(1'b1), .IN5(~na1866_1), .IN6(~na2763_1), .IN7(na79_1),
                      .IN8(na80_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6462_2 ( .OUT(na6462_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6462_1_i) );
// C_MX4b////      x104y65     80'h00_0018_00_0040_0AF7_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6463_1 ( .OUT(na6463_1), .IN1(na9947_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na9146_2), .IN5(~na9159_2), .IN6(~na9157_2), .IN7(~na82_1),
                      .IN8(na6673_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y64     80'h00_0018_00_0040_0A7F_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6464_1 ( .OUT(na6464_1), .IN1(na9947_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9146_2), .IN5(~na9156_2), .IN6(~na36_2), .IN7(~na82_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x112y47     80'h00_FE00_00_0040_0AE3_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6465_1 ( .OUT(na6465_1_i), .IN1(1'b1), .IN2(na67_2), .IN3(~na478_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na2763_1), .IN7(na6463_1),
                      .IN8(na6464_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6465_2 ( .OUT(na6465_1), .CLK(na4116_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6465_1_i) );
// C_MX4b////      x110y42     80'h00_0018_00_0040_0AFB_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6466_1 ( .OUT(na6466_1), .IN1(1'b1), .IN2(~na36_1), .IN3(na81_2), .IN4(1'b1), .IN5(~na1866_1), .IN6(~na9535_2), .IN7(na81_1),
                      .IN8(~na1865_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y108     80'h00_0018_00_0040_0A50_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6467_1 ( .OUT(na6467_1), .IN1(1'b1), .IN2(~na9168_2), .IN3(1'b1), .IN4(na9713_2), .IN5(na2703_1), .IN6(1'b0), .IN7(na1114_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y106     80'h00_0018_00_0040_0AC0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6468_1 ( .OUT(na6468_1), .IN1(1'b1), .IN2(na2919_1), .IN3(1'b1), .IN4(na92_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1033_1), .IN8(na9406_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y102     80'h00_0018_00_0040_0AC0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6469_1 ( .OUT(na6469_1), .IN1(1'b1), .IN2(na2919_1), .IN3(1'b1), .IN4(na92_1), .IN5(1'b0), .IN6(1'b0), .IN7(na9240_2), .IN8(na2705_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y102     80'h00_0018_00_0040_0A30_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6470_1 ( .OUT(na6470_1), .IN1(1'b1), .IN2(na2919_1), .IN3(1'b1), .IN4(~na92_1), .IN5(na2702_1), .IN6(na9407_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y104     80'h00_0018_00_0040_0A30_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6471_1 ( .OUT(na6471_1), .IN1(1'b1), .IN2(~na2919_1), .IN3(1'b1), .IN4(~na92_1), .IN5(na9408_2), .IN6(na892_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y106     80'h00_0018_00_0040_0A30_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6472_1 ( .OUT(na6472_1), .IN1(1'b1), .IN2(~na2919_1), .IN3(1'b1), .IN4(~na92_1), .IN5(na9409_2), .IN6(na2701_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x120y106     80'h00_0018_00_0040_0AC0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6473_1 ( .OUT(na6473_1), .IN1(1'b1), .IN2(~na2919_1), .IN3(1'b1), .IN4(na92_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1123_1), .IN8(na1079_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x124y98     80'h00_0018_00_0040_0A50_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6474_1 ( .OUT(na6474_1), .IN1(1'b1), .IN2(~na9168_2), .IN3(1'b1), .IN4(na9713_2), .IN5(na1342_1), .IN6(1'b0), .IN7(na2704_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y76     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6475_1 ( .OUT(na6475_1), .IN1(1'b1), .IN2(na1008_2), .IN3(1'b1), .IN4(na1009_1), .IN5(na4252_1), .IN6(na4261_1), .IN7(na1013_2),
                      .IN8(na4282_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y100     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6476_1 ( .OUT(na6476_1), .IN1(1'b1), .IN2(na980_1), .IN3(na2675_1), .IN4(1'b1), .IN5(na3214_2), .IN6(na5167_1), .IN7(na6066_1),
                      .IN8(na6078_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y58     80'h00_0018_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6477_1 ( .OUT(na6477_1), .IN1(1'b1), .IN2(~na1008_2), .IN3(1'b1), .IN4(na1009_1), .IN5(na4253_2), .IN6(na4244_1), .IN7(na4274_2),
                      .IN8(na236_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x122y58     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6478_1 ( .OUT(na6478_1), .IN1(1'b1), .IN2(~na1008_2), .IN3(1'b1), .IN4(~na1009_1), .IN5(na4275_1), .IN6(na239_2), .IN7(na4254_1),
                      .IN8(na4245_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x123y60     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6479_1 ( .OUT(na6479_1), .IN1(1'b1), .IN2(~na1008_2), .IN3(1'b1), .IN4(~na1009_1), .IN5(na4276_2), .IN6(na240_2), .IN7(na4255_2),
                      .IN8(na4246_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y59     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6480_1 ( .OUT(na6480_1), .IN1(1'b1), .IN2(na1008_2), .IN3(1'b1), .IN4(~na1009_1), .IN5(na241_2), .IN6(na4277_1), .IN7(na4247_2),
                      .IN8(na4256_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y60     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6481_1 ( .OUT(na6481_1), .IN1(1'b1), .IN2(~na1008_2), .IN3(1'b1), .IN4(~na1009_1), .IN5(na4278_2), .IN6(na242_2), .IN7(na4257_2),
                      .IN8(na4248_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y60     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6482_1 ( .OUT(na6482_1), .IN1(1'b1), .IN2(na1008_2), .IN3(1'b1), .IN4(~na1009_1), .IN5(na243_2), .IN6(na4279_2), .IN7(na4249_1),
                      .IN8(na4258_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x121y58     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6483_1 ( .OUT(na6483_1), .IN1(1'b1), .IN2(na1008_2), .IN3(1'b1), .IN4(na1009_1), .IN5(na4250_1), .IN6(na4259_2), .IN7(na244_2),
                      .IN8(na4280_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x119y55     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6484_1 ( .OUT(na6484_1), .IN1(1'b1), .IN2(na1008_2), .IN3(1'b1), .IN4(na1009_1), .IN5(na4251_2), .IN6(na4260_2), .IN7(na245_2),
                      .IN8(na4281_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x111y63     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6485_1 ( .OUT(na6485_1), .IN1(1'b1), .IN2(na3284_2), .IN3(1'b1), .IN4(~na1727_1), .IN5(na3285_1), .IN6(na5219_2), .IN7(na3282_1),
                      .IN8(na5215_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y114     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6486_1 ( .OUT(na6486_1), .IN1(1'b1), .IN2(~na980_1), .IN3(~na2675_1), .IN4(1'b1), .IN5(na6080_1), .IN6(na6068_1), .IN7(na5169_1),
                      .IN8(na107_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y114     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6487_1 ( .OUT(na6487_1), .IN1(1'b1), .IN2(~na980_1), .IN3(~na2675_1), .IN4(1'b1), .IN5(na6081_2), .IN6(na6069_2), .IN7(na5170_2),
                      .IN8(na116_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y117     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6488_1 ( .OUT(na6488_1), .IN1(1'b1), .IN2(na980_1), .IN3(na2675_1), .IN4(1'b1), .IN5(na3496_2), .IN6(na5171_1), .IN7(na6070_1),
                      .IN8(na6082_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x125y118     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6489_1 ( .OUT(na6489_1), .IN1(1'b1), .IN2(na980_1), .IN3(na2675_1), .IN4(1'b1), .IN5(na129_2), .IN6(na5172_2), .IN7(na6071_2),
                      .IN8(na6083_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y100     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6490_1 ( .OUT(na6490_1), .IN1(1'b1), .IN2(na980_1), .IN3(na2675_1), .IN4(1'b1), .IN5(na103_2), .IN6(na5178_2), .IN7(na6077_2),
                      .IN8(na6089_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x117y100     80'h00_0018_00_0040_0AF0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6491_1 ( .OUT(na6491_1), .IN1(1'b1), .IN2(na980_1), .IN3(~na2675_1), .IN4(1'b1), .IN5(na6074_1), .IN6(na6086_1), .IN7(na149_2),
                      .IN8(na5175_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x114y101     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6492_1 ( .OUT(na6492_1), .IN1(1'b1), .IN2(~na980_1), .IN3(~na2675_1), .IN4(1'b1), .IN5(na6088_1), .IN6(na6076_1), .IN7(na5177_1),
                      .IN8(na3499_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x118y100     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6493_1 ( .OUT(na6493_1), .IN1(1'b1), .IN2(na980_1), .IN3(na2675_1), .IN4(1'b1), .IN5(na3258_2), .IN6(na5176_2), .IN7(na6075_2),
                      .IN8(na6087_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x128y113     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6494_1 ( .OUT(na6494_1), .IN1(1'b1), .IN2(~na980_1), .IN3(na2675_1), .IN4(1'b1), .IN5(na5174_2), .IN6(na142_2), .IN7(na6085_2),
                      .IN8(na6073_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y118     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6495_1 ( .OUT(na6495_1), .IN1(1'b1), .IN2(na980_1), .IN3(na2675_1), .IN4(1'b1), .IN5(na3494_2), .IN6(na5168_2), .IN7(na6067_2),
                      .IN8(na6079_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x126y119     80'h00_0018_00_0040_0AF0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6496_1 ( .OUT(na6496_1), .IN1(1'b1), .IN2(na980_1), .IN3(~na2675_1), .IN4(1'b1), .IN5(na6072_1), .IN6(na6084_1), .IN7(na135_2),
                      .IN8(na5173_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x90y100     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6497_1 ( .OUT(na6497_1), .IN1(1'b1), .IN2(na3277_1), .IN3(na282_1), .IN4(1'b1), .IN5(na3287_2), .IN6(na5445_1), .IN7(na3278_2),
                      .IN8(na5449_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x81y88     80'h00_F600_00_0040_0AE0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6498_1 ( .OUT(na6498_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(1'b0), .IN6(na2594_1), .IN7(na2552_1),
                      .IN8(na5941_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6498_2 ( .OUT(na6498_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6498_1_i) );
// C_MX4b/D///      x77y75     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6499_1 ( .OUT(na6499_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5942_1), .IN6(na2553_1), .IN7(na2596_1),
                      .IN8(na3950_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6499_2 ( .OUT(na6499_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6499_1_i) );
// C_MX4b/D///      x57y85     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6500_1 ( .OUT(na6500_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5943_2), .IN6(na2554_1), .IN7(na2597_1),
                      .IN8(na9857_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6500_2 ( .OUT(na6500_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6500_1_i) );
// C_MX4b/D///      x80y82     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6501_1 ( .OUT(na6501_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5944_1), .IN6(na9614_2), .IN7(na2598_1),
                      .IN8(na3964_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6501_2 ( .OUT(na6501_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6501_1_i) );
// C_MX4b/D///      x77y81     80'h00_F600_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6502_1 ( .OUT(na6502_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na2599_1), .IN6(na9859_2), .IN7(na5945_2),
                      .IN8(na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6502_2 ( .OUT(na6502_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6502_1_i) );
// C_MX4b/D///      x78y81     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6503_1 ( .OUT(na6503_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5946_1), .IN6(na2557_1), .IN7(na2600_1),
                      .IN8(na3966_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6503_2 ( .OUT(na6503_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6503_1_i) );
// C_MX4b/D///      x78y89     80'h00_F600_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6504_1 ( .OUT(na6504_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na5830_2), .IN6(na9635_2), .IN7(na2558_1),
                      .IN8(na5947_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6504_2 ( .OUT(na6504_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6504_1_i) );
// C_MX4b/D///      x75y80     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6505_1 ( .OUT(na6505_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2559_1), .IN6(na5948_1), .IN7(na3968_1),
                      .IN8(na2602_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6505_2 ( .OUT(na6505_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6505_1_i) );
// C_MX4b/D///      x78y78     80'h00_F600_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6506_1 ( .OUT(na6506_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na5832_1), .IN6(na2603_1), .IN7(na2560_1),
                      .IN8(na5962_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6506_2 ( .OUT(na6506_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6506_1_i) );
// C_MX4b/D///      x74y80     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6507_1 ( .OUT(na6507_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5963_2), .IN6(na2561_1), .IN7(na2604_1),
                      .IN8(na3970_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6507_2 ( .OUT(na6507_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6507_1_i) );
// C_MX4b/D///      x79y87     80'h00_F600_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6508_1 ( .OUT(na6508_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na2605_1), .IN6(na5834_1), .IN7(na5964_2),
                      .IN8(na9620_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6508_2 ( .OUT(na6508_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6508_1_i) );
// C_MX4b/D///      x77y77     80'h00_F600_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6509_1 ( .OUT(na6509_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na2606_1), .IN6(na9854_2), .IN7(na5965_2),
                      .IN8(na2563_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6509_2 ( .OUT(na6509_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6509_1_i) );
// C_MX4b/D///      x73y91     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6510_1 ( .OUT(na6510_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na9621_2), .IN6(na5953_1), .IN7(na5836_2),
                      .IN8(na2607_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6510_2 ( .OUT(na6510_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6510_1_i) );
// C_MX4b/D///      x75y86     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6511_1 ( .OUT(na6511_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2565_1), .IN6(na5953_2), .IN7(na9855_2),
                      .IN8(na9638_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6511_2 ( .OUT(na6511_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6511_1_i) );
// C_MX4b/D///      x77y86     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6512_1 ( .OUT(na6512_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2566_1), .IN6(na9913_2), .IN7(na5838_1),
                      .IN8(na2609_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6512_2 ( .OUT(na6512_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6512_1_i) );
// C_MX4b/D///      x63y75     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6513_1 ( .OUT(na6513_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2574_2), .IN6(na5956_1), .IN7(na3945_1),
                      .IN8(na9640_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6513_2 ( .OUT(na6513_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6513_1_i) );
// C_MX4b/D///      x75y82     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6514_1 ( .OUT(na6514_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2576_2), .IN6(na5957_2), .IN7(na5840_1),
                      .IN8(na2611_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6514_2 ( .OUT(na6514_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6514_1_i) );
// C_MX4b/D///      x63y80     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6515_1 ( .OUT(na6515_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5958_1), .IN6(na2578_2), .IN7(na2612_1),
                      .IN8(na3947_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6515_2 ( .OUT(na6515_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6515_1_i) );
// C_MX4b/D///      x76y83     80'h00_F600_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6516_1 ( .OUT(na6516_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na9641_2), .IN6(na9910_2), .IN7(na9915_2),
                      .IN8(na2580_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6516_2 ( .OUT(na6516_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6516_1_i) );
// C_MX4b/D///      x69y80     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6517_1 ( .OUT(na6517_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na9631_2), .IN6(na5960_1), .IN7(na3949_1),
                      .IN8(na2614_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6517_2 ( .OUT(na6517_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6517_1_i) );
// C_MX4b/D///      x76y87     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6518_1 ( .OUT(na6518_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2584_2), .IN6(na9916_2), .IN7(na5844_2),
                      .IN8(na2615_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6518_2 ( .OUT(na6518_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6518_1_i) );
// C_MX4b/D///      x76y88     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6519_1 ( .OUT(na6519_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na9917_2), .IN6(na2586_2), .IN7(na2616_1),
                      .IN8(na3952_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6519_2 ( .OUT(na6519_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6519_1_i) );
// C_MX4b/D///      x80y90     80'h00_F600_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6520_1 ( .OUT(na6520_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na5846_2), .IN6(na2617_1), .IN7(na2588_2),
                      .IN8(na9919_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6520_2 ( .OUT(na6520_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6520_1_i) );
// C_MX4b/D///      x76y85     80'h00_F600_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6521_1 ( .OUT(na6521_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na2618_1), .IN6(na9856_2), .IN7(na5964_1),
                      .IN8(na2590_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6521_2 ( .OUT(na6521_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6521_1_i) );
// C_MX4b/D///      x79y86     80'h00_F600_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6522_1 ( .OUT(na6522_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na2619_1), .IN6(na5848_1), .IN7(na5965_1),
                      .IN8(na2592_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6522_2 ( .OUT(na6522_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6522_1_i) );
// C_MX4b/D///      x78y85     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6523_1 ( .OUT(na6523_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5967_2), .IN6(na2567_1), .IN7(na2620_1),
                      .IN8(na3956_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6523_2 ( .OUT(na6523_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6523_1_i) );
// C_MX4b/D///      x79y88     80'h00_F600_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6524_1 ( .OUT(na6524_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na5850_2), .IN6(na2621_1), .IN7(na2568_1),
                      .IN8(na9924_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6524_2 ( .OUT(na6524_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6524_1_i) );
// C_MX4b/D///      x78y90     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6525_1 ( .OUT(na6525_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2569_1), .IN6(na9929_2), .IN7(na3958_1),
                      .IN8(na9644_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6525_2 ( .OUT(na6525_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6525_1_i) );
// C_MX4b/D///      x78y92     80'h00_F600_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6526_1 ( .OUT(na6526_1_i), .IN1(1'b1), .IN2(~na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na2570_1), .IN6(na9927_2), .IN7(na5852_1),
                      .IN8(na9645_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6526_2 ( .OUT(na6526_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6526_1_i) );
// C_MX4b/D///      x79y89     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6527_1 ( .OUT(na6527_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5971_2), .IN6(na2571_1), .IN7(na2624_1),
                      .IN8(na3960_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6527_2 ( .OUT(na6527_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6527_1_i) );
// C_MX4b/D///      x80y92     80'h00_F600_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6528_1 ( .OUT(na6528_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(~na42_2), .IN5(na2625_1), .IN6(na5854_1), .IN7(na9930_2),
                      .IN8(na2572_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6528_2 ( .OUT(na6528_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6528_1_i) );
// C_MX4b/D///      x75y84     80'h00_F600_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6529_1 ( .OUT(na6529_1_i), .IN1(1'b1), .IN2(na45_1), .IN3(1'b1), .IN4(na42_2), .IN5(na5972_1), .IN6(na9628_2), .IN7(na9646_2),
                      .IN8(na9858_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6529_2 ( .OUT(na6529_1), .CLK(na4116_1), .EN(~na3243_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6529_1_i) );
// C_MX4b////      x68y83     80'h00_0018_00_0040_0AB0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6530_1 ( .OUT(na6530_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na356_1), .IN6(na3280_1), .IN7(1'b0), .IN8(na9595_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x68y81     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6531_1 ( .OUT(na6531_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2595_1), .IN6(na9596_2), .IN7(na354_1),
                      .IN8(na3359_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y79     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6532_1 ( .OUT(na6532_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2391_1), .IN6(na2393_1), .IN7(na2423_1),
                      .IN8(na3361_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y76     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6533_1 ( .OUT(na6533_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2392_1), .IN6(na2394_1), .IN7(na2424_1),
                      .IN8(na3363_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y82     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6534_1 ( .OUT(na6534_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na9597_2), .IN6(na2393_1), .IN7(na3365_2),
                      .IN8(na2425_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y84     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6535_1 ( .OUT(na6535_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2396_1), .IN6(na2394_1), .IN7(na3367_1),
                      .IN8(na2426_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y84     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6536_1 ( .OUT(na6536_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na2427_1), .IN6(na3369_2), .IN7(na2395_1),
                      .IN8(na2397_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y82     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6537_1 ( .OUT(na6537_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2396_1), .IN6(na9598_2), .IN7(na2428_1),
                      .IN8(na3371_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y83     80'h00_0018_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6538_1 ( .OUT(na6538_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na3373_1), .IN6(na2429_1), .IN7(na2399_1),
                      .IN8(na2397_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y84     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6539_1 ( .OUT(na6539_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na2430_1), .IN6(na3375_2), .IN7(na2398_1),
                      .IN8(na9599_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y84     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6540_1 ( .OUT(na6540_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na2431_1), .IN6(na3377_1), .IN7(na2399_1),
                      .IN8(na2401_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y86     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6541_1 ( .OUT(na6541_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na2432_1), .IN6(na3379_2), .IN7(na2400_1),
                      .IN8(na2402_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y86     80'h00_0018_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6542_1 ( .OUT(na6542_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na3381_2), .IN6(na2433_1), .IN7(na2403_1),
                      .IN8(na2401_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y88     80'h00_0018_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6543_1 ( .OUT(na6543_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na3383_1), .IN6(na2434_1), .IN7(na2404_1),
                      .IN8(na2402_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y87     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6544_1 ( .OUT(na6544_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na2435_1), .IN6(na3385_2), .IN7(na2403_1),
                      .IN8(na2405_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y80     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6545_1 ( .OUT(na6545_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na2436_1), .IN6(na3387_1), .IN7(na2404_1),
                      .IN8(na2406_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y86     80'h00_0018_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6546_1 ( .OUT(na6546_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na3389_1), .IN6(na2437_1), .IN7(na2407_1),
                      .IN8(na2405_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y89     80'h00_0018_00_0040_0AF0_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6547_1 ( .OUT(na6547_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na3391_2), .IN6(na2438_1), .IN7(na2408_1),
                      .IN8(na2406_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y88     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6548_1 ( .OUT(na6548_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2409_1), .IN6(na9600_2), .IN7(na3393_1),
                      .IN8(na2439_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y90     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6549_1 ( .OUT(na6549_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na9601_2), .IN6(na2410_1), .IN7(na9609_2),
                      .IN8(na3395_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x54y91     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6550_1 ( .OUT(na6550_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2409_1), .IN6(na2411_1), .IN7(na2441_1),
                      .IN8(na3397_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y90     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6551_1 ( .OUT(na6551_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2412_1), .IN6(na2410_1), .IN7(na3399_1),
                      .IN8(na9611_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y92     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6552_1 ( .OUT(na6552_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2413_1), .IN6(na2411_1), .IN7(na3401_1),
                      .IN8(na9612_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y86     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6553_1 ( .OUT(na6553_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2412_1), .IN6(na2414_1), .IN7(na2444_1),
                      .IN8(na3403_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y90     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6554_1 ( .OUT(na6554_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2413_1), .IN6(na2415_1), .IN7(na2445_1),
                      .IN8(na3405_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y92     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6555_1 ( .OUT(na6555_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2416_1), .IN6(na2414_1), .IN7(na3407_2),
                      .IN8(na2446_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y93     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6556_1 ( .OUT(na6556_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2417_1), .IN6(na2415_1), .IN7(na3409_2),
                      .IN8(na2447_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y92     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6557_1 ( .OUT(na6557_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2416_1), .IN6(na2418_1), .IN7(na2448_1),
                      .IN8(na3411_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x58y91     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6558_1 ( .OUT(na6558_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2417_1), .IN6(na9602_2), .IN7(na2449_1),
                      .IN8(na3413_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y92     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6559_1 ( .OUT(na6559_1), .IN1(1'b1), .IN2(~na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2420_1), .IN6(na2418_1), .IN7(na3415_1),
                      .IN8(na2450_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y90     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6560_1 ( .OUT(na6560_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(na48_1), .IN5(na2451_1), .IN6(na3417_2), .IN7(na2419_1),
                      .IN8(na2421_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y86     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6561_1 ( .OUT(na6561_1), .IN1(1'b1), .IN2(na55_1), .IN3(1'b1), .IN4(~na48_1), .IN5(na2420_1), .IN6(na3332_1), .IN7(na2390_1),
                      .IN8(na3419_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x76y123     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a6562_2 ( .OUT(na6562_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a6562_6 ( .COUTY1(na6562_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6562_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x135y110     80'h00_0078_00_0020_0C66_C5CF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a6563_1 ( .OUT(na6563_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na8394_1), .IN6(1'b1), .IN7(1'b1), .IN8(na4079_1),
                      .CINX(1'b0), .CINY1(na6624_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a6563_4 ( .OUT(na6563_2), .COUTY1(na6563_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4079_2), .IN5(~na8394_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na4079_1), .CINX(1'b0), .CINY1(na6624_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x135y111     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a6565_1 ( .OUT(na6565_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na4081_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na6563_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a6565_4 ( .OUT(na6565_2), .COUTY1(na6565_4), .IN1(1'b1), .IN2(1'b1), .IN3(na4081_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4081_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na6563_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x135y112     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a6567_1 ( .OUT(na6567_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na4083_1),
                      .CINX(1'b0), .CINY1(na6565_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a6567_4 ( .OUT(na6567_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4083_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na4083_1),
                      .CINX(1'b0), .CINY1(na6565_4), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a6569 ( .Y(na6569_1), .I(cdone_ice40) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a6570 ( .Y(na6570_1), .I(clk10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6571 ( .O(core_en_ice40), .A(na8423_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6572 ( .Y(na6572_1), .O(creset_ice40), .A(na8424_10), .EN(na8425_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6573 ( .Y(na6573_1), .O(gatemate_debug_3), .A(na8426_10), .EN(na8427_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6574 ( .Y(na6574_1), .O(gatemate_debug_4), .A(na8428_10), .EN(na8429_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6575 ( .Y(na6575_1), .O(gatemate_debug_5), .A(na8430_10), .EN(na8431_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6576 ( .O(hyperram_clk_n), .A(na8432_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6577 ( .O(hyperram_clk_p), .A(na8433_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6578 ( .O(hyperram_cs_n), .A(na8434_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6579 ( .Y(na6579_1), .O(hyperram_dq[0]), .A(na8435_10), .EN(na8436_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6580 ( .Y(na6580_1), .O(hyperram_dq[1]), .A(na8437_10), .EN(na8438_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6581 ( .Y(na6581_1), .O(hyperram_dq[2]), .A(na8439_10), .EN(na8440_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6582 ( .Y(na6582_1), .O(hyperram_dq[3]), .A(na8441_10), .EN(na8442_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6583 ( .Y(na6583_1), .O(hyperram_dq[4]), .A(na8443_10), .EN(na8444_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6584 ( .Y(na6584_1), .O(hyperram_dq[5]), .A(na8445_10), .EN(na8446_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6585 ( .Y(na6585_1), .O(hyperram_dq[6]), .A(na8447_10), .EN(na8448_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6586 ( .Y(na6586_1), .O(hyperram_dq[7]), .A(na8449_10), .EN(na8450_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6587 ( .O(hyperram_rst_n), .A(na8451_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6588 ( .Y(na6588_1), .O(hyperram_rwds), .A(na8452_10), .EN(na8453_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6589 ( .Y(_d7), .O(i2c0_scl), .A(na8454_10), .EN(na8455_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6590 ( .Y(na6590_1), .O(i2c0_sda), .A(na8456_10), .EN(na8457_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6591 ( .Y(_d8), .O(i2c1_scl), .A(na8458_10), .EN(na8459_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6592 ( .Y(na6592_1), .O(i2c1_sda), .A(na8460_10), .EN(na8461_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6593 ( .Y(na6593_1), .O(ice40_io_vcore_0), .A(na8462_10), .EN(na8463_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6594 ( .Y(na6594_1), .O(ice40_io_vcore_1), .A(na8464_10), .EN(na8465_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6595 ( .Y(na6595_1), .O(ice40_io_vcore_2), .A(na8466_10), .EN(na8467_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6596 ( .Y(na6596_1), .O(ice40_io_vcore_4), .A(na8468_10), .EN(na8469_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6597 ( .Y(na6597_1), .O(ice40_io_vio_0), .A(na8470_10), .EN(na8471_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6598 ( .Y(na6598_1), .O(ice40_io_vio_1), .A(na8472_10), .EN(na8473_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6599 ( .Y(na6599_1), .O(ice40_io_vio_2), .A(na8474_10), .EN(na8475_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6600 ( .Y(na6600_1), .O(ice40_io_vio_3), .A(na8476_10), .EN(na8477_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6601 ( .Y(na6601_1), .O(ice40_io_vio_4), .A(na8478_10), .EN(na8479_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a6602 ( .Y(na6602_1), .O(ice40_io_vio_5), .A(na8480_10), .EN(na8481_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6603 ( .O(osc_en_ice40), .A(na8482_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a6604 ( .Y(na6604_1), .I(power_fauld_ice40) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6605 ( .O(spi_flash_clk), .A(na8483_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6606 ( .O(spi_flash_cs_n), .A(na8484_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a6607 ( .Y(na6607_1), .I(spi_flash_miso) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6608 ( .O(spi_flash_mosi), .A(na8485_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6609 ( .O(spi_ice40_clk), .A(na8486_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6610 ( .O(spi_ice40_cs_n), .A(na8487_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a6611 ( .Y(na6611_1), .I(spi_ice40_miso) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6612 ( .O(spi_ice40_mosi), .A(na8488_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a6613 ( .Y(na6613_1), .I(uart_ice40_rx) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6614 ( .O(uart_ice40_tx), .A(na8489_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a6615 ( .Y(na6615_1), .I(uart_logging_rx) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6616 ( .O(uart_logging_tx), .A(na8490_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a6617 ( .Y(na6617_1), .I(usb_uart_rx) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6618 ( .O(usb_uart_tx), .A(na8491_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6619 ( .O(user_led_n0), .A(na8492_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6620 ( .O(user_led_n1), .A(na8493_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6621 ( .O(user_led_n2), .A(na8494_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6622 ( .O(user_led_n3), .A(na8495_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a6623 ( .O(vio_en_ice40), .A(na8496_10) );
// C_/C_0_1///      x135y109     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a6624_2 ( .OUT(na6624_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a6624_6 ( .COUTY1(na6624_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6624_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND/DST//AND/DST      x108y86     80'h20_BE00_80_0000_0C88_CF00
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6626_1 ( .OUT(na6626_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na6626_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0000)) 
           _a6626_2 ( .OUT(na6626_1), .CLK(na4116_1), .EN(1'b1), .SR(na3334_2), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6626_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6626_4 ( .OUT(na6626_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0100)) 
           _a6626_5 ( .OUT(na6626_2), .CLK(na4116_1), .EN(1'b1), .SR(na3334_2), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na6626_2_i) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_19_08_08_28_82),
             .REF_CLK(10.00),
             .OUT_CLK(8.00),
             .LOW_JITTER(1),
             .CI_FILTER_CONST(2),
             .CP_FILTER_CONST(4)) 
           _a6627 ( .USR_PLL_LOCKED_STDY(_d9), .USR_PLL_LOCKED(na6627_2), .CLK270(na6627_3), .CLK180(na6627_4), .CLK90(na6627_5), .CLK0(na6627_6),
                    .CLK_REF_OUT(_d10), .CLK_REF(na6662_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
CC_USR_RSTN            _a6628 ( .USR_RSTN(na6628_1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_00_00_C0_00_1B_00_00_23_03_13_23_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6629 ( .DOA({_d11, _d12, _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23, _d24, _d25, _d26, _d27, _d28,
                   _d29, _d30, na6629_21, na6629_22, na6629_23, na6629_24, na6629_25, na6629_26, na6629_27, na6629_28, na6629_29, na6629_30,
                   na6629_31, na6629_32, na6629_33, na6629_34, na6629_35, na6629_36, na6629_37, na6629_38, na6629_39, na6629_40}),
                    .DOAX({_d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44, _d45, _d46, _d47, _d48,
                   _d49, _d50, _d51, _d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65, _d66, _d67,
                   _d68, _d69, _d70}),
                    .DOB({_d71, _d72, _d73, _d74, _d75, _d76, _d77, _d78, _d79, _d80, _d81, _d82, _d83, _d84, _d85, _d86, _d87, _d88,
                   _d89, _d90, _d91, _d92, _d93, _d94, _d95, _d96, _d97, _d98, na6629_109, na6629_110, na6629_111, na6629_112, na6629_113,
                   na6629_114, na6629_115, na6629_116, na6629_117, na6629_118, na6629_119, na6629_120}),
                    .DOBX({_d99, _d100, _d101, _d102, _d103, _d104, _d105, _d106, _d107, _d108, _d109, _d110, _d111, _d112, _d113, _d114,
                   _d115, _d116, _d117, _d118, _d119, _d120, _d121, _d122, _d123, _d124, _d125, _d126, _d127, _d128, _d129, _d130, _d131,
                   _d132, _d133, _d134, _d135, _d136, _d137, _d138}),
                    .ECC1B_ERRA({_d139, _d140, _d141, _d142}),
                    .ECC1B_ERRB({_d143, _d144, _d145, _d146}),
                    .ECC2B_ERRA({_d147, _d148, _d149, _d150}),
                    .ECC2B_ERRB({_d151, _d152, _d153, _d154}),
                    .FORW_CAS_WRAO(_d155), .FORW_CAS_WRBO(_d156), .FORW_CAS_BMAO(_d157), .FORW_CAS_BMBO(_d158), .FORW_CAS_RDAO(_d159),
                    .FORW_CAS_RDBO(_d160), .FORW_UADDRAO({_d161, _d162, _d163, _d164, _d165, _d166, _d167, _d168, _d169, _d170, _d171,
                   _d172, _d173, _d174, _d175, _d176}),
                    .FORW_LADDRAO({_d177, _d178, _d179, _d180, _d181, _d182, _d183, _d184, _d185, _d186, _d187, _d188, _d189, _d190,
                   _d191, _d192}),
                    .FORW_UADDRBO({_d193, _d194, _d195, _d196, _d197, _d198, _d199, _d200, _d201, _d202, _d203, _d204, _d205, _d206,
                   _d207, _d208}),
                    .FORW_LADDRBO({_d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216, _d217, _d218, _d219, _d220, _d221, _d222,
                   _d223, _d224}),
                    .FORW_UA0CLKO(_d225), .FORW_UA0ENO(_d226), .FORW_UA0WEO(_d227), .FORW_LA0CLKO(_d228), .FORW_LA0ENO(_d229), .FORW_LA0WEO(_d230),
                    .FORW_UA1CLKO(_d231), .FORW_UA1ENO(_d232), .FORW_UA1WEO(_d233), .FORW_LA1CLKO(_d234), .FORW_LA1ENO(_d235), .FORW_LA1WEO(_d236),
                    .FORW_UB0CLKO(_d237), .FORW_UB0ENO(_d238), .FORW_UB0WEO(_d239), .FORW_LB0CLKO(_d240), .FORW_LB0ENO(_d241), .FORW_LB0WEO(_d242),
                    .FORW_UB1CLKO(_d243), .FORW_UB1ENO(_d244), .FORW_UB1WEO(_d245), .FORW_LB1CLKO(_d246), .FORW_LB1ENO(_d247), .FORW_LB1WEO(_d248),
                    .CLOCKA({_d249, _d250, _d251, _d252}),
                    .CLOCKB({_d253, _d254, _d255, _d256}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, na6646_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na6649_10, na6652_9, na6654_10, na6656_9, na6658_10, na6660_9, na6667_10, na6669_9, na6670_10, na6676_9,
                   na6679_10, na6680_9, na6682_10, na6683_9, na6685_10, na6686_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({na6687_10, na6688_9, na6689_10, na6690_9, na6691_10, na6693_9, na6694_10, na6697_9, na6698_10, na6703_9,
                   na6704_10, na6707_9, na6708_10, na6713_9, na6714_10, na6715_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na6716_10, na6717_9, na6718_10, na6720_9, na6721_10, na6722_9, na6725_10, na6726_9, na6728_10, na6729_9,
                   na6730_10, na6731_9, na6732_10, na6734_9, na6735_10, na6737_9, na6738_10, na6739_9, na6740_10, na6742_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na6744_10, na6746_9, na6747_10, na6748_9, na6751_10,
                   na6754_9, na6755_10, na6756_9, na6757_10, na6758_9, na6760_10, na6761_9}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na6762_10, na6763_9, na6764_10, na6765_9, na6766_10, na6772_9, na6773_10, na6785_9, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_00_06_00_00_C3_03_13_23_00_00_23_00_13_23_00_00_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6630 ( .DOA({na6630_1, na6630_2, na6630_3, na6630_4, na6630_5, na6630_6, na6630_7, na6630_8, na6630_9, na6630_10, na6630_11,
                   na6630_12, na6630_13, na6630_14, na6630_15, na6630_16, na6630_17, na6630_18, na6630_19, na6630_20, _d257, _d258,
                   _d259, _d260, _d261, _d262, _d263, _d264, _d265, _d266, _d267, _d268, _d269, _d270, _d271, _d272, _d273, _d274, _d275,
                   _d276}),
                    .DOAX({_d277, _d278, _d279, _d280, _d281, _d282, _d283, _d284, _d285, _d286, _d287, _d288, _d289, _d290, _d291,
                   _d292, _d293, _d294, _d295, _d296, _d297, _d298, _d299, _d300, _d301, _d302, _d303, _d304, _d305, _d306, _d307, _d308,
                   _d309, _d310, _d311, _d312, _d313, _d314, _d315, _d316}),
                    .DOB({_d317, _d318, _d319, _d320, _d321, _d322, _d323, _d324, na6630_89, na6630_90, na6630_91, na6630_92, na6630_93,
                   na6630_94, na6630_95, na6630_96, na6630_97, na6630_98, na6630_99, na6630_100, _d325, _d326, _d327, _d328, _d329,
                   _d330, _d331, _d332, _d333, _d334, _d335, _d336, _d337, _d338, _d339, _d340, _d341, _d342, _d343, _d344}),
                    .DOBX({_d345, _d346, _d347, _d348, _d349, _d350, _d351, _d352, _d353, _d354, _d355, _d356, _d357, _d358, _d359,
                   _d360, _d361, _d362, _d363, _d364, _d365, _d366, _d367, _d368, _d369, _d370, _d371, _d372, _d373, _d374, _d375, _d376,
                   _d377, _d378, _d379, _d380, _d381, _d382, _d383, _d384}),
                    .ECC1B_ERRA({_d385, _d386, _d387, _d388}),
                    .ECC1B_ERRB({_d389, _d390, _d391, _d392}),
                    .ECC2B_ERRA({_d393, _d394, _d395, _d396}),
                    .ECC2B_ERRB({_d397, _d398, _d399, _d400}),
                    .FORW_CAS_WRAO(_d401), .FORW_CAS_WRBO(_d402), .FORW_CAS_BMAO(_d403), .FORW_CAS_BMBO(_d404), .FORW_CAS_RDAO(_d405),
                    .FORW_CAS_RDBO(_d406), .FORW_UADDRAO({_d407, _d408, _d409, _d410, _d411, _d412, _d413, _d414, _d415, _d416, _d417,
                   _d418, _d419, _d420, _d421, _d422}),
                    .FORW_LADDRAO({_d423, _d424, _d425, _d426, _d427, _d428, _d429, _d430, _d431, _d432, _d433, _d434, _d435, _d436,
                   _d437, _d438}),
                    .FORW_UADDRBO({_d439, _d440, _d441, _d442, _d443, _d444, _d445, _d446, _d447, _d448, _d449, _d450, _d451, _d452,
                   _d453, _d454}),
                    .FORW_LADDRBO({_d455, _d456, _d457, _d458, _d459, _d460, _d461, _d462, _d463, _d464, _d465, _d466, _d467, _d468,
                   _d469, _d470}),
                    .FORW_UA0CLKO(_d471), .FORW_UA0ENO(_d472), .FORW_UA0WEO(_d473), .FORW_LA0CLKO(_d474), .FORW_LA0ENO(_d475), .FORW_LA0WEO(_d476),
                    .FORW_UA1CLKO(_d477), .FORW_UA1ENO(_d478), .FORW_UA1WEO(_d479), .FORW_LA1CLKO(_d480), .FORW_LA1ENO(_d481), .FORW_LA1WEO(_d482),
                    .FORW_UB0CLKO(_d483), .FORW_UB0ENO(_d484), .FORW_UB0WEO(_d485), .FORW_LB0CLKO(_d486), .FORW_LB0ENO(_d487), .FORW_LB0WEO(_d488),
                    .FORW_UB1CLKO(_d489), .FORW_UB1ENO(_d490), .FORW_UB1WEO(_d491), .FORW_LB1CLKO(_d492), .FORW_LB1ENO(_d493), .FORW_LB1WEO(_d494),
                    .CLOCKA({_d495, _d496, _d497, _d498}),
                    .CLOCKB({_d499, _d500, _d501, _d502}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na6791_10, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1({na6793_10, na6795_9, na6800_10, na6801_9, na6802_10, na6804_9, na6806_10, na6808_9, na6809_10, na6811_9,
                   na6813_10, na6814_9, na6815_10, na6817_9, na6818_10, na6819_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({na6820_10, na6821_9, na6822_10, na6824_9, na6825_10, na6826_9, na6827_10, na6829_9, na6830_10, na6831_9,
                   na6832_10, na6833_9, na6835_10, na6837_9, na6838_10, na6840_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na6842_10, na6843_9, na6844_10, na6846_9, na6848_10, na6850_9, na6851_10, na6852_9, na6854_10, na6856_9, na6857_10,
                   na6858_9, na6860_10, na6861_9, na6862_10, na6863_9, na6865_10, na6872_9, na6873_10, na6874_9, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na6876_10, na6877_9, na6878_10, na6880_9, na6882_10, na6883_9,
                   na6884_10, na6885_9, na6890_10, na6893_9, na6894_10, na6895_9, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({na6897_10, na6898_9, na6899_10, na6901_9, na6902_10, na6903_9, na6905_10, na6906_9, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'hbceef9cc631cef3bcef39de779cc6318c6318c6318c6318df318c6318c6318c6318c639ce739ce6f),
             .INIT_01(320'h9be739be739be739be739de6318c6318c6318e6798e6f1dc6399e7318c631ccf33cdef9ceef98c73),
             .INIT_02(320'hbce777ce6f9cdf3bcef3bce777ce6f9cdf37ceef9be737cdf3bcef3bce777ce6f9cdf37ce737cdf3),
             .INIT_03(320'h9ceef9ce73bce739be739ce737ce739ce6f9ce739cdf39be739be739ce739be739cdf39cdf3bcef3),
             .INIT_04(320'h7cef3bcef39dc631cdf39ce73bce73b8e6f9ce73bbe6f9ce73bbe739ce779be739ce779ce771be73),
             .INIT_05(320'h18c739dc639be739ceef7ce739cef39be739ceef7ce739cef39be739cee71ce7798e737ce739dc63),
             .INIT_06(320'h1cdf39ce777be739ce779ce777ce739de739cef39ddf39ce739de739de737ce739dc639cee31ce77),
             .INIT_07(320'h9ce73b8e739ce739cc739be739cef398e737ce739dc739ce739ce639cdf39ce779cc739be739cee3),
             .INIT_08(320'h9ce73bce6f9ce73bcdf39ce73bce6f9ce73bbdf39ce73bcc631ce739ce7398e737ce739de731ce6f),
             .INIT_09(320'h9de73bbe739ce73b8c739be739cee39ce739ce731ce6f9ce73bce639cdf39ce7718e6f9ce73bbdf3),
             .INIT_0A(320'h9ce73bce639cdf39ce7798e737ce739dc779cc737ce739dc7398eef7ce739cef39ceef9ce73bce73),
             .INIT_0B(320'h7be779de779cef398ee3b8c771de7398e737ce739de731ce6f9ce73bcc739be739cee3bce731ce6f),
             .INIT_0C(320'hbbdf39ce63b8e771ddef9ce731dc73b8ee39dc777be739cc771cee3b8c777cef3bcef39de731dc77),
             .INIT_0D(320'h9cef39be739ceef7ce739cef39be739cee3b8e7718c6398df39ce731de7398de31cdf39dc771cee3),
             .INIT_0E(320'h9cdf39ce779cc737ce739dc63bbe779de779cee3bbe779de779cee3bbe779de779cee3bbc777ce73),
             .INIT_0F(320'h7ce739cef39be739cee398ee3b8de3bbe739ce779cdf39ce771cc6f9de779de73b8c739ce739ce63),
             .INIT_10(320'h7ce739cc739be739cef31dc7718eef9de779de73bcc731dc777be779de779cef31cc771dc63bbc77),
             .INIT_11(320'h9ce777be739ce779cdf39ce771dc63b8ee318c7318e731dc7798ee31ce639be739ceef1bc7798ee3),
             .INIT_12(320'h1ce6f9ce73b8e731ce6f9ce73bce639cdf39ce7798e737ce739dc731cdf39ce777be739ce779cdf3),
             .INIT_13(320'h1ce631be779de779cee31bdf3bcef3bce7718c637be739ce779cdf39ce771dc639cc739be739cef3),
             .INIT_14(320'hbbe739cef39ce779ceef9cc739ce779cc739be739ceef98c639cc739ce739ce739ce739ce7398e73),
             .INIT_15(320'h18e6f9be739ce779ce777ce739de739cef39ddf39ce739de731cc639cdf39ce777cdf39ce73bce73),
             .INIT_16(320'h3ce739ce739ce7398e7398c7399e739ce739ce739cc739cc639ccf398c6318c6318c6318c73b8c63),
             .INIT_17(320'h98c6398c7318c7318de318c631cc6398c6398c6f18e739ce739ce739ce739ce7398e731ce631cc73),
             .INIT_18(320'h98c6399e7318c733cc739cc6318c7318c731cc6378e6398e731ce631bc7398e7318de398e631ce63),
             .INIT_19(320'h1be63b8c739ce7318c6318c6318c631ce639ce639cc731ce7318e6398e639cc6318e679ce631ccf3),
             .INIT_1A(320'h98e731ce771ce6f9ce6f9ce7398c6318e731ce731ce6398e737ce739cc6318c631cc6398c6398c6f),
             .INIT_1B(320'h1ce6398e7718e731ce731ce639cee39ce739ce6318c7398e7398e731cc739be739ce6318c7398e73),
             .INIT_1C(320'h9ce639dc73b8c7398e7398e731ce771ce731ce7398e771cee31cdf39ce739ce7318c631ce639ce63),
             .INIT_1D(320'h18c6318c6318e6798e6f9ce6318e777cc6318c6318c631ccf318e731ce639ce639cc739dc739cc73),
             .INIT_1E(320'h18c639cc6318c6318c631be7398c639ddf318c6318c6318c733cc7318c6318c637ce7318c73bbe63),
             .INIT_1F(320'h18e6799e679cc631ccf31cc6318c6318c6318df39cc6f9ce6318e777cc6318c6318c631ccf31cc63),
             .INIT_20(320'h9cc631ce6398e631be7318c6318e679cc639cc6398ee378e771bc7318c6318e679cc631ccf398c63),
             .INIT_21(320'h98c631ccf31cde39cc631cc637ce6318c733cc737cdf39cc6318e6798e6f9be7398c631ccf31cde3),
             .INIT_22(320'h3ccf33cc7398e6f1cc6399e739ce6318c733cc7378df398c6378c7318e6798e739be7318de378df3),
             .INIT_23(320'h18c6318c6318c6318c733cc7378e7718e6798e6f1cee31ccf31ce6f9dc733ce6318e679cc6318c73),
             .INIT_24(320'h1be779de779ceef9de779de73b8c6399e639cc73b8c731be7398e6318e6378c6399e639be639dc63),
             .INIT_25(320'h9de73bbc737ce6378df3bcef3bce777ce6378e6f9cc6f9bc6f9be731bc6f9de779de73bbe639dc63),
             .INIT_26(320'h1ccf31cdf3bcef3bce777be779de779cee318e6f98e779be6398e7318e6f18c737ce6f9ce6f9de77),
             .INIT_27(320'h18c6318c6318e6799e6798e739cde31ccf31cdf318e6798e6f98c733cc7398c631cc6f9ce6378c63),
             .INIT_28(320'h18e6f9ce7318c6318e6798e737cef3bcef39dc637cc731be631cdf39ce6318df318c631cc6399e73),
             .INIT_29(320'h98c639be739ce739ce6398c637be739ce731cc631bdf39ce739ce731cc631bc73b8e639dc73b8c63),
             .INIT_2A(320'hb8e6f9cdf31de7378c771cdf39cdf318e6f98c6318e6318e6798e739cc6f9de779de73b8c737ce73),
             .INIT_2B(320'h18c6318e631ccf33ccf318e6f9ce7398e6318c739cc739de631ce7798df3bcef3bce771cdf39bc63),
             .INIT_2C(320'h9de73bce739bc7318c739ce6f1be779de779cee318e637cc639be7398c637cc6318e679cc6318c63),
             .INIT_2D(320'h9ce73bce6f18c733cc739be7398c6318e6798e737cc779be7378c6399e631ce6f1cc6398c6f9de77),
             .INIT_2E(320'h7ce7318c631ccf31cdf39cc6318c7318e6798e6f9ce6318c6398c733cc737ce7318c631cc6399e63),
             .INIT_2F(320'h3ce6318c6318c631ccf33ccf31cdf39cc6318c7318e6798e739cdf39cc6318e739bc7318e6798e73),
             .INIT_30(320'h3cc737cdf39ce7318c631ccf31ce6f9de779de73b8c6f98e637cc639be739cc631be6318c6398c73),
             .INIT_31(320'h98c737ce7398c6318c6318e6798e6f1be7398e6318c739ce739cee39ce7398c737ce7398c6318c73),
             .INIT_32(320'h18c6318c739ce7398e739ce631ce739ce639ce7398c739ce739cee39ce7398c739ce739cee39ce73),
             .INIT_33(320'h18c739ce7398e739ce631ce739ce639ce7398c737ce7398c6318c6399e639be7398e6318c6318c63),
             .INIT_34(320'h7cc779cdf31de6f98df37cc779cdf31de6f98de398c731cc631cdf39ce6318c6399e639be7398e63),
             .INIT_35(320'h98de398c731cc631cdf39ce6318c6399e639cdf39ce6318c6399e639cdf37cc779cdf31de6f98df3),
             .INIT_36(320'h9cdf39ce6318c6399e639cdf37cc779cdf31de6f98df37cc779cdf31de6f98df37cc779cdf31de6f),
             .INIT_37(320'h1de6f98df37cc779cdf31de6f98df37cc779cdf31de6f98de398c731cc631cdf39ce6318c6399e63),
             .INIT_38(320'h9cdf31de6f98de398c731cc631cdf39ce6318c6399e639cdf39ce6318c6399e639cdf37cc779cdf3),
             .INIT_39(320'h18c6399e639cdf39ce6318c6399e639cdf37cc779cdf31de6f98df37cc779cdf31de6f98df37cc77),
             .INIT_3A(320'h9cdf31de737cc7378c63bbc63b8e6318c6318c6398c6398c6398c6398c731ce639cc731be739ce63),
             .INIT_3B(320'h7cc7378c63bbc63b8e6318c6318c6398c6398c6398c6398c731ce639cc731be739ce6318c6399e63),
             .INIT_3C(320'h1cc6398e6318e639cc7398e637ce739cc6318e639cc7398e637ce739cc6318c6399e639cdf31de73),
             .INIT_3D(320'h9be739bc7378df37cc779cdf31de6f9ce737ce6f9ce6f1cde37cdf31de737cc779cdf39cde39bc6f),
             .INIT_3E(320'h9cc731be739ce6318c731ce639cc731be739ce6318c631ccf318e737cdf31de737cc779be739cdf3),
             .INIT_3F(320'h9be739ce739ce739be737ce7378e6f1be6f98ef39be63bce6f9ce6f1cde378e631cc7318c731ce63),
             .INIT_40(320'h1cee31dc6f1cc6318c6399e6799e631ce6f9be63bcdf39ce739ce739cdf39be739bc7378df37cc77),
             .INIT_41(320'h18c731bc731cc6f1cde39cdf31ce6398de398e6398c733cc7378c6399e639bc6378e639dc639dc6f),
             .INIT_42(320'h3cc7378e6f1cde398c733cc731bc6318e6378e6398e7318c6398de39bc7378e6318e6798e631cde3),
             .INIT_43(320'h1ce631ccf31cc6f18e6f1bc7398de378de398de39cc6f18e639cc6399e639bc7378e6f1cde398c73),
             .INIT_44(320'h1bc731bc7398de31cc7318e6318e6798e6378c731ce6f18e7378de39cc6f1bc6f1cc6f1ce6378c73),
             .INIT_45(320'h98e7318e6798e739cde39ce7398e7398c731ce631ccf318e6f18c631cc639bc7318de378e731bc6f),
             .INIT_46(320'h3cc7378de39ce7398de39cc6f1cc6f1ce6378c731cc7398c733cc7378de398de398de39cc6f18e63),
             .INIT_47(320'h9cc631bc7378e631ccf31cde39bc7378e6f1cc6399e6398c631cc6318e737cc7778e631cee318c73),
             .INIT_48(320'h18c6378e6318c631ccf31cdf318e6398c6318de398c6318de398c6318c733cc739be631bc7378e63),
             .INIT_49(320'h18c631ccf33ccf31cdf318e6398c6318de398c6318de398c6318c733cc737cc6398e6318c6378e63),
             .INIT_4A(320'h1cc6399e639be7398c631ccf31cdf39cc6318e679ce63b8de39dc6f1cc6318c631ccf398c6399e73),
             .INIT_4B(320'h98c6318c6f18c6399e639cdf398c6f9ce6318c733cc7378e6318c6399e639bc7398c6318e6798e6f),
             .INIT_4C(320'h99e7398c733ce631ce679ce6f98c6399e7318c733ce6318c6399e6799e7318c733cc739cc7318c6f),
             .INIT_4D(320'h9cc73b8e6f1bc739be6f18e6798e731cc63b8de398c73b8de398c6318c6f9ce7398c631ccf398c73),
             .INIT_4E(320'h9ce6318c739cee31be631ccf318e7318c731ce7398c639cc631cc7398c737ce631bc631ce639dc63),
             .INIT_4F(320'h1cc6399e639be7398c737ce6318c733cc737cdf39ce631cdef9cee31be7398c6f9ce6318c63bcc77),
             .INIT_50(320'h18c7378e6318e6798e7318c6398de398e631bc6318c733cc7398e739cdf398c737ce7318df398c63),
             .INIT_51(320'h99e6398c639cc6318e6398c639dc771cdf31cee3b8e6f18ef31de6f18c733cc7318c7398c631cc73),
             .INIT_52(320'h99e639cc7398e6f18e6378e6398c6f18c6399e739ce6318c6399e739cc6398c6f98c7318c6318c63),
             .INIT_53(320'h1ce737ce6318e739be7318c739cdf398c637ce6318c733cc7378e737cc7398c7318e6318c6318c63),
             .INIT_54(320'h98e6f9de779de73bbc7398e6f98c7798e631cdf31dc63b8c733ce631dc733ccf33cc7378e7718c63),
             .INIT_55(320'h18e6798e6f9ce63bbe73b8c631ce737ce639cc6398c7318ee318c6318c6399e7318ee318e6799e67),
             .INIT_56(320'h7cc6f18df398df318c6399e7318c6318c6399e6799e639be7398eef98e7318e631cc63b8c6318c63),
             .INIT_57(320'h9cc6f98c6318c6399e631cdf318c631cc639be7318c6f1bc637ce637cc6318c631ccf31cc6f98c73),
             .INIT_58(320'h7cc6398e739be631cc739cdf318e6f98df398df318c733cc639be6318c6398c737ce6318de378c6f),
             .INIT_59(320'h99e639bc6f98df398c6f18df398df31bc639bc731cc631ccf31cdf31be731be731be6318e6798e63),
             .INIT_5A(320'h18c739ce631bc6318c6399e639bc6f98c6318e637ce6398c6378de31be731be6378c7378e6318c63),
             .INIT_5B(320'h78e6318e6798e6f1be6378c6f9cc6f98de31cde398c6399e639cc6318e631bc731cc6398c6398c73),
             .INIT_5C(320'h1be731be6318e6798e6f1be6378c6f9cc6f98de31cde398c6399e639bc6f98de31be731be6378c73),
             .INIT_5D(320'h7cc6f9cc6f98c6399e639be7398c6f9ce7318df39ce6318c6399e639be637ce637cc631ccf31cdf3),
             .INIT_5E(320'hbce7778e7778e779ce6f9de779de73bbe779de779cee398c6399e639ce739bc631ccf31cc6f98c73),
             .INIT_5F(320'h18e637cef31ce6378df3bbe779de779ceef1cef39cdf3bcef3bce7778e779de6f1cef39cdf3bcef3),
             .INIT_60(320'h1be771cc6398c6318e731be7798e731bc6f9ddf3b8e631cc631cc7398df3bcc7398de37ceef9dc73),
             .INIT_61(320'h7be779de779cee318c631ccf398e6799e6798c731be779de779cef39cde39cde37be779de779cee3),
             .INIT_62(320'h98c637cdf378e631cc7318c6399e6318e6318df318c631ccf31be779de779cee319e6318c6318c63),
             .INIT_63(320'h9cee318e6798e6f1dc6399e639bc7718e6798e6f1dc6399e7318c631ccf33ccf31ce6f98c6798c63),
             .INIT_64(320'h3cc7378e6f1cde39be7398e637ce7398e637ce7398e637ce6398df39cc731be731cc6f9ce7798df3),
             .INIT_65(320'h99e639be631cc6399e639be631cc6399e639be731be731be731be7398df39cc6f9ce637ce7318c73),
             .INIT_66(320'h18c6318e6799e679cc639cc7318e739ce639ce779cc6398e739cc739cc6f1cc6399e639be631cc63),
             .INIT_67(320'h98c7318e631cc631cc6318c639be6318c7318c7318c639be6318c6f98e739be6318e7718c733ce63),
             .INIT_68(320'h9ce7318c737ce6f9be739ce7398e771cef318df39ce6318e6f9cdf37ce631cc631ccf31ce639bc73),
             .INIT_69(320'hbce739cef39ceef9ce739ce771ce73bce739dc739ce771ce73bcc739cef79dc6399e631cdf398c6f),
             .INIT_6A(320'h9ce739ce771ce73bce739dc739cee39ce7798e739def3b8c733cc639de6f1ce739de739ceef9ce73),
             .INIT_6B(320'h9ce7318e733ce739cc639ccf39ce7318e733cc639de6f1ce739de739ceef9ce73bce739cef39ceef),
             .INIT_6C(320'h1ce6318c731cc6378c6318c7318e6318e631bc639ce739ce739ce739ce739ce639cc7398c731ccf3),
             .INIT_6D(320'h1ce6398de39ce6318c6318e6798e7398c6318e6318e631bc731cc7398c6f1ce6318e6398c7318c73),
             .INIT_6E(320'h98c6318c6318c6318c631ce639ce639cc731ce739ce7318c639cc739cc7398e639ce739ce739cc73),
             .INIT_6F(320'h18c631ce7398c631cc6398c6398e6378c739ce6318df31ce739cc6318e731ce731ce6398e739ce73),
             .INIT_70(320'h9cc731ce6f9ce7398c631ce639ce639cc731ce739ce739ce639cdf39ce7318c639cc739be739ce63),
             .INIT_71(320'h18c637cc639ce7318c639cc739cc7398e639cdf39ce7318c639be739be739ce6318e631ce639ce63),
             .INIT_72(320'h99e739ce731cee39dc6399e739ce7318c6399e6318e7318c637cc7318e631be639ce639cdf39ce73),
             .INIT_73(320'h3ccf31cdf3bcef3bce7718e6f9cc6f9cc6f9de779de73bbc6399e6398ee37ce6398df398c6399e67),
             .INIT_74(320'h18e6798e739be639ce771be6398c6399e639bde398e739dc6398c631ccf398c6399e7318c631ccf3),
             .INIT_75(320'h7ce7398df39ce6318e6799e6798e6f9cc739cee398c6f98e739dc631ccf31cdef1cc739cee31cc63),
             .INIT_76(320'h7ce731be7398c6318c6318e771be739cc6318c6318c6318c6f9ce7318e6318c637ce7398df39ce63),
             .INIT_77(320'h1bc639ce6318e7318c631be73b8c6f9cc637ce631be7318df39cc637ce7798c6f9ce737ce737ce63),
             .INIT_78(320'h98e637cef3bcef39dc7318de39cc6f18c6318e7318c631ccf31ce6f9de779de73b8e739be631be63),
             .INIT_79(320'hbce771cc631ce737cc6378c739de6f9cc6f9de779de73b8e631be6398df3bcef3bce771cc6378e73),
             .INIT_7A(320'h98c6318c6f9de779de73b8e631bc7318e631cc6398c7318e637cef3bcef39dc7318c7378df3bcef3),
             .INIT_7B(320'h1ce731cde39cc6398de31ce6318e7398e6f1ce631cc6398c6f9de779de73b8e631bde39bde39ce63),
             .INIT_7C(320'h18de398c631ce731cde39cc6398de31ce6318e7398e6f1ce631cc6398c6f9de779de73b8e631bc63),
             .INIT_7D(320'hb8e6318e7318df3bcef3bce771cc631cdf31ce7378c7398c639cc639bc737bc737cef3bcef39dc73),
             .INIT_7E(320'h78df3bcef3bce7718df3bcef3bce771cdf31cce31cc631cc6378de39ce6398de39cc6f9de779de73),
             .INIT_7F(320'h18df3bcef3bce771cc637cc639cc637cef3bcef39dc7318df318c631cc6f9de779de73bcc7318c63)) 
           _a6631 ( .DOA({_d503, _d504, _d505, _d506, _d507, _d508, _d509, _d510, _d511, _d512, _d513, _d514, _d515, _d516, _d517, _d518,
                   _d519, _d520, _d521, _d522, _d523, _d524, _d525, _d526, _d527, _d528, _d529, _d530, _d531, _d532, _d533, _d534, _d535,
                   _d536, _d537, na6631_36, na6631_37, na6631_38, na6631_39, na6631_40}),
                    .DOAX({_d538, _d539, _d540, _d541, _d542, _d543, _d544, _d545, _d546, _d547, _d548, _d549, _d550, _d551, _d552,
                   _d553, _d554, _d555, _d556, _d557, _d558, _d559, _d560, _d561, _d562, _d563, _d564, _d565, _d566, _d567, _d568, _d569,
                   _d570, _d571, _d572, _d573, _d574, _d575, _d576, _d577}),
                    .DOB({_d578, _d579, _d580, _d581, _d582, _d583, _d584, _d585, _d586, _d587, _d588, _d589, _d590, _d591, _d592, _d593,
                   _d594, _d595, _d596, _d597, _d598, _d599, _d600, _d601, _d602, _d603, _d604, _d605, _d606, _d607, _d608, _d609, _d610,
                   _d611, _d612, _d613, _d614, _d615, _d616, _d617}),
                    .DOBX({_d618, _d619, _d620, _d621, _d622, _d623, _d624, _d625, _d626, _d627, _d628, _d629, _d630, _d631, _d632,
                   _d633, _d634, _d635, _d636, _d637, _d638, _d639, _d640, _d641, _d642, _d643, _d644, _d645, _d646, _d647, _d648, _d649,
                   _d650, _d651, _d652, _d653, _d654, _d655, _d656, _d657}),
                    .ECC1B_ERRA({_d658, _d659, _d660, _d661}),
                    .ECC1B_ERRB({_d662, _d663, _d664, _d665}),
                    .ECC2B_ERRA({_d666, _d667, _d668, _d669}),
                    .ECC2B_ERRB({_d670, _d671, _d672, _d673}),
                    .FORW_CAS_WRAO(_d674), .FORW_CAS_WRBO(_d675), .FORW_CAS_BMAO(_d676), .FORW_CAS_BMBO(_d677), .FORW_CAS_RDAO(_d678),
                    .FORW_CAS_RDBO(_d679), .FORW_UADDRAO({_d680, _d681, _d682, _d683, _d684, _d685, _d686, _d687, _d688, _d689, _d690,
                   _d691, _d692, _d693, _d694, _d695}),
                    .FORW_LADDRAO({_d696, _d697, _d698, _d699, _d700, _d701, _d702, _d703, _d704, _d705, _d706, _d707, _d708, _d709,
                   _d710, _d711}),
                    .FORW_UADDRBO({_d712, _d713, _d714, _d715, _d716, _d717, _d718, _d719, _d720, _d721, _d722, _d723, _d724, _d725,
                   _d726, _d727}),
                    .FORW_LADDRBO({_d728, _d729, _d730, _d731, _d732, _d733, _d734, _d735, _d736, _d737, _d738, _d739, _d740, _d741,
                   _d742, _d743}),
                    .FORW_UA0CLKO(_d744), .FORW_UA0ENO(_d745), .FORW_UA0WEO(_d746), .FORW_LA0CLKO(_d747), .FORW_LA0ENO(_d748), .FORW_LA0WEO(_d749),
                    .FORW_UA1CLKO(_d750), .FORW_UA1ENO(_d751), .FORW_UA1WEO(_d752), .FORW_LA1CLKO(_d753), .FORW_LA1ENO(_d754), .FORW_LA1WEO(_d755),
                    .FORW_UB0CLKO(_d756), .FORW_UB0ENO(_d757), .FORW_UB0WEO(_d758), .FORW_LB0CLKO(_d759), .FORW_LB0ENO(_d760), .FORW_LB0WEO(_d761),
                    .FORW_UB1CLKO(_d762), .FORW_UB1ENO(_d763), .FORW_UB1WEO(_d764), .FORW_LB1CLKO(_d765), .FORW_LB1ENO(_d766), .FORW_LB1WEO(_d767),
                    .CLOCKA({_d768, _d769, _d770, _d771}),
                    .CLOCKB({_d772, _d773, _d774, _d775}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na6907_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na6908_10, na6910_9, na6911_10, na6912_9, na6914_10, na6915_9, na6916_10, na6918_9, na6919_10, na6920_9,
                   na6922_10, na6923_9, na6924_10, na6926_9, na6927_10, na6928_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na6930_10, na6931_9, na6932_10, na6934_9, na6939_10,
                   na6940_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h62103820341c20c62103421081a398a4080e629062398a10e80c4310c4310c4310c4310000000003),
             .INIT_01(320'he1d0ce1d0ce1d0ce1d09a54110c4310c4310c503410074363140d000e3818a060180671a1234046c),
             .INIT_02(320'hed31d3a387470e8eb3b0ed31d3a387470e83a3a741d1c3a0e8eb3b0ed31d3a387470e83a19c3a0e8),
             .INIT_03(320'he73a74779ceb214c1d1c642983a38c8530747190a60e8e1d0ce1d0c8731ca1d0c870e8670e8eb3b0),
             .INIT_04(320'h3a3acec3b4c767caf0e86779cee79cee7874779ce9d074779ce9d0cef39dc1d0cef39dcf39de9d1d),
             .INIT_05(320'h4b79de763ce1d1de73a33a19de73b8e1d1de73a33a19de73b8e1d1de73a3e779dc5f1c3a3bce74fc),
             .INIT_06(320'he70e8ef39d19d0cef39dcf39d3a190e7698ce33de74f0a713ce773ce759c3a3bce74b8ef3a1c779d),
             .INIT_07(320'h4779cec79cef39ce739ce1d1de73a42739c3a3bce773ce779ce739ce70e8ef39d2139ce1d1de73a5),
             .INIT_08(320'h6779cee3874779ce80e86779cee3874779ce8ce86779cee07c4f39de739ce739c3a3bce7484e7387),
             .INIT_09(320'hc67bce9e14e279ced30ce1d1de73a9e73bce739ce73874779ce909ce70e8ef39d8f3874779ce8ce8),
             .INIT_0A(320'h4779ce979ce70e8ef39d2739c3a3bce743dc779c3a3bce747ce73a33a19de73b9e73a74321ced319),
             .INIT_0B(320'h19d0963611a633c073b8e8f9d8f71de739c3a3bce74bce73874779ce939ce1d1de73b1ee3bce7387),
             .INIT_0C(320'he8ce867398ecf9dc74674339cc767cee3a3e771d19d0ce731d9f3b8e8f9d3a12c6c234c6780e771d),
             .INIT_0D(320'he73b8e1d1de73a33a19de73b8e1d1de73a1e871dbe391e70e867399e773ce6071af0e86771d9f3b8),
             .INIT_0E(320'he70e8ef39d2139c3a3bce767ce9d0963611a633ce9d0963611a633ce9d0963611a633ce8c3d3a19d),
             .INIT_0F(320'h3a19de73b8e1d1de73b3ef3b4ee061e9d0cef39dc70e8ef39d9f3074258d84698cf33ce779ce739c),
             .INIT_10(320'h3a190e7298e1d1de73a5e771d1f3a74258d84698c831de771d19d0963611a6320c779dc767ce8c3d),
             .INIT_11(320'hef39d19d0cef39dc70e8ef39d0f67cee3b7c703ce07bd84431673b4c779cc1d1de73a308c3dcf3b8),
             .INIT_12(320'he73874779cec7bce73874779ce979ce70e8ef39d2739c3a3bce74bde70e8ef39d19d0cef39dc70e8),
             .INIT_13(320'he1383e1d0963611a633c00ce84b1b08d319e007c19d0cef39dc70e8ef39d9f701ef39ce1d1de73a4),
             .INIT_14(320'he9d0c873b4c6719ef3a78531c4f39dc638ce1d1de73a743214e703ce279ce42b4c10086b31cc4718),
             .INIT_15(320'h0c50301d0cef39dcf39d3a190e7698ce33de74f0a713ce7694e6798670e8ef39d1a0e86779cee79c),
             .INIT_16(320'h1a11ce739de739ce7318e733c40d08e739cef39ce7398c7399e20680071c8e381c7238e0798ec431),
             .INIT_17(320'hef303e607cc379de60710df1c8f381ef298ef3038c79c4f39ce63bca1010ad11cc05086418988228),
             .INIT_18(320'h4739140d08e72281a00842387c723ce071dc77981879c0071dc73bcc0c38ee39de6073c0f1c0e3b8),
             .INIT_19(320'h88f93ee13ce73bce6391c71b8e271c2e694c6301ac214e631ce2785e278de62310c5034239c8a068),
             .INIT_1A(320'hc56b0853bda6387433874739de731c01734a63180d610a731c3a39cef398e5f1c8f395ef298ef303),
             .INIT_1B(320'h2e694c63bdc0734a6318ed610a77b4c639ce779cc70b9a5318c06b085398e1d1ce779cc7339a5318),
             .INIT_1C(320'he779ced719cf039a5318c76b0853bda631dc739de73b5c673c0f0e86739ce73bce63944e694c6318),
             .INIT_1D(320'h8531c886218c503410074339c0f31d3a190a63910c4318a0680111c4e694c6305ac214ef698c771c),
             .INIT_1E(320'h0f221c5381e4781e4781e1d0ce703cc74e864298e44310c6281a0808f1bc4f03c3a19ce0798e9d0c),
             .INIT_1F(320'h0c50300c034003c8a0682003c8f03c0f23c0f0e8673874339c0f31d3a190a63910c4318a0682003c),
             .INIT_20(320'h6739c0f79ccf31c89d1ce72218c5034023cc739c0073c18719e0e781f23c0c5034239c8a0680071c),
             .INIT_21(320'h673918a068200e86739c0f3913a39ce46281a0803a0e86739c8c5034100741d0ce73918a068200e8),
             .INIT_22(320'h180601a08005f874023140d08e779ce72281a0803a0e8673983a1bc8c5034111ce1d1ce70e83a0e8),
             .INIT_23(320'hc0698e4701a63910c6281a0803a19d8c50341007433b18a06822387476281a11ce450340038e0628),
             .INIT_24(320'hc1d1d6761da63a74759d87698e863140d04002fcee23ce1d0ce73bcc729c1c63140d0401d01c6791),
             .INIT_25(320'h87698e9d0c3a39c3a0e8eb3b0ed31d3a39c3a1874738741d0741d1ce1d074759d87698e9d0ca761c),
             .INIT_26(320'h8a068200e8eb3b0ed31d19d1d6761da63a3e5f83e4f9dc1d0ce4f9ce37874363c3a387433874759d),
             .INIT_27(320'h0e2340d31c0c50300c034111cef0f18a068200e88c50341007446281a08001f988f3874339c1c431),
             .INIT_28(320'he67874321ce73018c5034111c3a12c6c234c679c1f27cc1d1cef0e86439ce60e8e471c6f23140d00),
             .INIT_29(320'he739801d10a739ce739c6739819d0c85294a739cc0ce88539ce739ce339cc0c78ccf03c6678cf038),
             .INIT_2A(320'he8787470e86771c3a19d8f0e8670e8e70074707ce27910c5034111ce73874258d84698cf23c3a190),
             .INIT_2B(320'ha0698e77818a060180680100743214a539ce603de7399e771c0f79dc70e84b1b08d319070e8e1d0c),
             .INIT_2C(320'h84698cf004e1d00e707cef38741d0963611a633ce4f983a39de1d0c873983a3910c50340238e0711),
             .INIT_2D(320'h473bdee387446281a088e1d0c873988c5034111c3a19dc1d1c3a23140d002238743391e72274258d),
             .INIT_2E(320'h3a190e73118a068200e86429ce613c8c5034100743214e7309e46281a0803a190a73984f23140d04),
             .INIT_2F(320'h1a001c4681a63818a06018068200e86429ce613c8c5034111ce70e86439cc5f9ce1d008c5034111c),
             .INIT_30(320'h1a0803a0e86429ce73118a068223874258d84698cf383e4f983a39de1d0c8739cc1d1c8e38de4628),
             .INIT_31(320'he733c3a190e7398886218c5034100741d0c8539ce633ce779cef3b4c639ce733c3a190e73980c628),
             .INIT_32(320'h0e381c733ce779ce7318e739ccf39de739cc639ce733ce779cef3b4c639ce733ce779cef3b4c639c),
             .INIT_33(320'he63bce779ce7318e739cef39de739cc639ce73bc3a190e73988863140d0401d0c8539ce6238e471c),
             .INIT_34(320'h3a19dc70e8677074707c3a19dc70e86770747063c0e789e39ccf0e86439ce623140d0401d0c8539c),
             .INIT_35(320'h47063c0e789e39ccf0e86439ce623140d04470e86439ce623140d044707c3a19dc70e8677074707c),
             .INIT_36(320'h470e86439ce623140d044707c3a19dc70e8677074707c3a19dc70e8677074707c3a19dc70e867707),
             .INIT_37(320'h677074707c3a19dc70e8677074707c3a19dc70e86770747063c0e789e39ccf0e86439ce623140d04),
             .INIT_38(320'hc70e86770747063c0e789e39ccf0e86439ce623140d04470e86439ce623140d044707c3a19dc70e8),
             .INIT_39(320'he223140d04470e86439ce623140d044707c3a19dc70e8677074707c3a19dc70e8677074707c3a19d),
             .INIT_3A(320'h470e86771c3a19c3a23ce8e3cecf98e4f9c1f383e6393e6393e6381e703dc779ccf398e1d90a639c),
             .INIT_3B(320'h3a19c3a23ce8e3cecf98e4f9c1f383e6393e6393e6381e703dc779ccf398e1d90a639ce223140d04),
             .INIT_3C(320'h9e063c0f1ce07b8ef399e731c3b214c739c447b8ef399e731c3b214c739c4443140d04470e86771c),
             .INIT_3D(320'he1d0ce1d003a07c3a19dc70e8677074739c3a38743387400e81f0e86771c3a19dc70e8670e801d03),
             .INIT_3E(320'hcf398e1d90a639ce223dc779ccf398e1d90a639ce22218a0680111c1f0e86771c3a19dc1d1ce70e8),
             .INIT_3F(320'hc1d1cef3bce639ce1d1c3a19c3a00740f87433b8e1d0cee38743387400e81cf031e278e703dc779c),
             .INIT_40(320'h0e33c8e7831e07c8863140c0300d0022383e1d0cee0e8e779de731ce70e8e1d0ce1d003a07c3a19d),
             .INIT_41(320'hbf03ce1d0cef387430e86707c9f3bcc7061e778de46281a0803a23140d0401d0c3a001c6791c6783),
             .INIT_42(320'h1a0803a187430e8646281a088e1d17e079c3a19dee39ce739de70e860c3c3a19d8c5034111cef0e8),
             .INIT_43(320'h6e3918a068223874778741d0c870e83a0e8670e8643874278dc723140d0401d0c3a187430e864628),
             .INIT_44(320'h41d0ce1d0c870e80f13c6c7910c5034111c3a33de63874679c3a0e86438741d07433874321c3a13c),
             .INIT_45(320'he371c8c5034111cef0e86739cef318e713c6e3918a0680100741f98cf381e1d01c70793a190e1d07),
             .INIT_46(320'h1a0803a0e86739ce70e867387433874321c3a03c4f1b8e46281a0803a0e8670e8670e86438741789),
             .INIT_47(320'he739ce1d0c3a1918a068200e861d0c3a1874323140d0400781e639c0f31c3a19d1871c9f3b80c628),
             .INIT_48(320'he639c18f989f0318a068200e8e7001c7398e7061c7398e7063e627c0c6281a088e0f93e1d0c3a19d),
             .INIT_49(320'h0e3818a06018068200e8e7001c7398e7061c7398e7063e627c0c6281a0803a39c0071ce639c1871c),
             .INIT_4A(320'h4323140d0401d0ce73918a068200e86739c8c50340011cf071c67839e07c0e3818a0684739140d00),
             .INIT_4B(320'hef313e62274063140d04470e8e73874339ce46281a0803a19ce063140d0401d0ce73818c50341007),
             .INIT_4C(320'h40d001f2281a11c8fd03400631cf9140d08e72281a001c703140c0300d08e72281a088e7799e6383),
             .INIT_4D(320'hef398e878740e3de1c070c503410008e381cf071c7038cf063c0f85e078743218e70318a0684723f),
             .INIT_4E(320'hc771ce071de633ce1d118a068010003f23de639dc703cc739c0f798a73983a39ce1d11e779cc767c),
             .INIT_4F(320'h6f23140d0401d0ce73983a39ce46281a0803a0e8ef71ce50e7433b8e1d0ce73874339ce6381ee79d),
             .INIT_50(320'he72fc3a01d8c503410003f311e70e8673bcc0e310c6281a08005f9ce70e8e73803a19ce70e867398),
             .INIT_51(320'h40d04470bcc739cef3bcc7383e771d3f07c9f3b8e8f87447b8e7403ec6281a088e1798e739de7798),
             .INIT_52(320'h40d04000fcef3074479c3a19cef3038863140d08e73bce639140d08e779cc7383ef398e707ce6391),
             .INIT_53(320'h8f39c3a39ce579ce1d1ce733ce70e8e739d3a39ce46281a0803a19c3a190e623ce47910c43108631),
             .INIT_54(320'h410074759d87698e8efcef3074339d0079c8f0e8e747cec6281a011c7628180601a0803a18de6290),
             .INIT_55(320'h8c503410074331ce9d908d31c0111c3a190a7311e703c1f3b10c6218863140d000e3a3e450300c03),
             .INIT_56(320'h3a387430e8670e8e063140d008e034c703140c0300d0401d0cc73a74321cc479c0f07cec4310c431),
             .INIT_57(320'h43387470310c43140d00200e8e5f988f381e1d01e628389d0c3a19c3a381886218a06822387473bc),
             .INIT_58(320'h3a391ef31ce1d1c8f798e70e8e4787470e8670e8e46281a00401d1cbf311e703c3a03cc50713a187),
             .INIT_59(320'h40d0401d07470e866387430e8670e8e1d17e1d00ef0318a068200e8e1d0ce1d0ce1d1c8c5034111c),
             .INIT_5A(320'he603dc73bcc0e218863140d0401d07472fcc479c3a19cef3141c4e861d0ce1d1c3a2fc3a00188631),
             .INIT_5B(320'h3a0018c5034100741d1c3a18743387470e8bf0e80063140d04000fcc47bcc1d10a77986f311e0f99),
             .INIT_5C(320'he1d0ce1d1c8c5034100741d1c3a18743387470e8bf0e80063140d0401d07470e861d0ce1d1c3a2fc),
             .INIT_5D(320'h3a387433874723140d0401d0cc63874339ce60e86739cc063140d0401d1c3a19c3a3918a068200e8),
             .INIT_5E(320'hed31d3a19d3a19d853874759d87698e9d1d6761da63bde443140d04473bce1d118a06822387473bc),
             .INIT_5F(320'hc679c3a3ace779c1e4e8e9d1d6761da63a7433b0a70e8eb3b0ed31d3a19d87687433b0a70e8eb3b0),
             .INIT_60(320'he1d1d3f311e73a3c73bce1d1d673bce0e27474e8e9f98af39d1f31de70e8eb39de70753a3a7476fc),
             .INIT_61(320'h19d0963611a633c9f0318a0680450300c0340088e1d0963611a633c070e8070e819d1d6761da63a3),
             .INIT_62(320'he739c1f07c18f031e278e723cc1d18c739ce707c9f3918a06821d1d6761da63b1e1d18c739ce071c),
             .INIT_63(320'h643b88c503410074363140d0401d0d8c503410074363140d000e3818a0601806822383e07874631c),
             .INIT_64(320'h1a0803a187430e861d0c8639c3a190e731c3a190e731c3a198e70e867398e1d0cc73874321dc70e8),
             .INIT_65(320'h40d0401d1c6f23140d0401d1c6f23140d0401d1ce1d1ce1d1ce1d0ce70e8673874339c3a19ce4628),
             .INIT_66(320'he071c0c50300c0342397e7438e679cef39cef295e7791a721ce7398c7383cf03140d0401d1c6f231),
             .INIT_67(320'h87398e5f988f691a439cc6795e1d1ce663da4690e731de1d1ce4783e4f9ce1d1ce471d0c6281a011),
             .INIT_68(320'h43218e723c3a38741d10e739dc6339e77aca70e86431ce6787470e83a19ce02218a06822381e1d0c),
             .INIT_69(320'hed319ad33dce3a785389ad39d676b4ee738e7438ee71d6f6b4ee23dce03d4d43140d00200e867387),
             .INIT_6A(320'h85389ad39d676b4ee738e743dce3aded69dc47b9c07a9a86281a0044d407433b5a7739c73a74321c),
             .INIT_6B(320'h4739ce67881a11ce7399e20684739ce67881a0044d407433b5a7739c73a74321ced319ad33dce3a7),
             .INIT_6C(320'hc73bcc379dc77981e437c723ce07bca63bcc0e31e713ce7398ef284042b44730142190626208a068),
             .INIT_6D(320'he631ce70e86739c886310c50340108472fcc679c0e3b8e0c3ce0038ee3830e3b8e4f13c707cc279d),
             .INIT_6E(320'he731caf31c8f31c6f31c6e694c6309ac214e631ce73bce6389cd298c60b58429cc639cef39ce739c),
             .INIT_6F(320'hc7007c739de731ccf399ed31cce39c1e47ce779cc707c9f318ef398e1734a63180d610a7318e739d),
             .INIT_70(320'hac214e63874739de731cee694c6319ac214e631ce779ce739cef0e8e73bce63840039de1d1ce779c),
             .INIT_71(320'he63801f278e73bce6389cd298c60b58429cc70e8e73bce6391e1d0ce1d1ce779cc701c4e694c6305),
             .INIT_72(320'h00d08e73bce76b8ce79140d08e73bce639140d040111c0f31c1f27ce731ce0f93e779cef0e8e73bc),
             .INIT_73(320'h18068200e84b1b08d319e478747387473874759d87698e9e3140d040073c3a198e70e86723140c03),
             .INIT_74(320'h8c50341100e1d1cef319e0f93e623140d0400ce8673bcc6793e60318a0684739140d000e3818a060),
             .INIT_75(320'h3a190e70e86439c8c50300c03410074339de633ca7227473bcc67918a068200674339de633c9f301),
             .INIT_76(320'h3a19ce1d0ce72218871483319e1d0c87391e078de6795e47874321ce071caf23c3a190e70e86439c),
             .INIT_77(320'he0e3cc639ce071dc639ce1d0cee3874339c3a19ce1d0ce70e86739c3a19dc73874321c3a19c3a39c),
             .INIT_78(320'he731c3a3acec3b4c767cc70e86738745799e4f9ce72218a068223874759d87698edf9ce1d1ce1d1c),
             .INIT_79(320'hed31d9f31c9f39c3a39c18799e7707473874759d87698ecf98e0f91c70e8eb3b0ed31d9f31c3a190),
             .INIT_7A(320'hc707ce63874759d87698ecf98e0e7cc4f989f313e627cc4f983a3acec3b4c767cc703c3a0e8eb3b0),
             .INIT_7B(320'h0f79cc50e86039cc7071e639ce07bce62874301ce6383e63874759d87698ecf98e0ce860ce86439c),
             .INIT_7C(320'hc7075c72bc0f79cc50e86039cc7075e639ce07bce62874301ce6383e63874759d87698ecf98e0e3c),
             .INIT_7D(320'hecf98e0f98e70e8eb3b0ed31d9f31cbf07c9f39c3a27ce7383e739c01d0c19d0c3a3acec3b4c767c),
             .INIT_7E(320'h1e4e84b1b08d319e70e8eb3b0ed31d9f07c9f0e8e739c9f31c3a0e86439cc70e8673874759d87698),
             .INIT_7F(320'he70e8eb3b0ed31d1f31c1f1bcc739c3a3acec3b4c767cc707cbe39ccf3874258d84698cf39de639c)) 
           _a6632 ( .DOA({_d776, _d777, _d778, _d779, _d780, _d781, _d782, _d783, _d784, _d785, _d786, _d787, _d788, _d789, _d790, _d791,
                   _d792, _d793, _d794, _d795, _d796, _d797, _d798, _d799, _d800, _d801, _d802, _d803, _d804, _d805, _d806, _d807, _d808,
                   _d809, _d810, na6632_36, na6632_37, na6632_38, na6632_39, na6632_40}),
                    .DOAX({_d811, _d812, _d813, _d814, _d815, _d816, _d817, _d818, _d819, _d820, _d821, _d822, _d823, _d824, _d825,
                   _d826, _d827, _d828, _d829, _d830, _d831, _d832, _d833, _d834, _d835, _d836, _d837, _d838, _d839, _d840, _d841, _d842,
                   _d843, _d844, _d845, _d846, _d847, _d848, _d849, _d850}),
                    .DOB({_d851, _d852, _d853, _d854, _d855, _d856, _d857, _d858, _d859, _d860, _d861, _d862, _d863, _d864, _d865, _d866,
                   _d867, _d868, _d869, _d870, _d871, _d872, _d873, _d874, _d875, _d876, _d877, _d878, _d879, _d880, _d881, _d882, _d883,
                   _d884, _d885, _d886, _d887, _d888, _d889, _d890}),
                    .DOBX({_d891, _d892, _d893, _d894, _d895, _d896, _d897, _d898, _d899, _d900, _d901, _d902, _d903, _d904, _d905,
                   _d906, _d907, _d908, _d909, _d910, _d911, _d912, _d913, _d914, _d915, _d916, _d917, _d918, _d919, _d920, _d921, _d922,
                   _d923, _d924, _d925, _d926, _d927, _d928, _d929, _d930}),
                    .ECC1B_ERRA({_d931, _d932, _d933, _d934}),
                    .ECC1B_ERRB({_d935, _d936, _d937, _d938}),
                    .ECC2B_ERRA({_d939, _d940, _d941, _d942}),
                    .ECC2B_ERRB({_d943, _d944, _d945, _d946}),
                    .FORW_CAS_WRAO(_d947), .FORW_CAS_WRBO(_d948), .FORW_CAS_BMAO(_d949), .FORW_CAS_BMBO(_d950), .FORW_CAS_RDAO(_d951),
                    .FORW_CAS_RDBO(_d952), .FORW_UADDRAO({_d953, _d954, _d955, _d956, _d957, _d958, _d959, _d960, _d961, _d962, _d963,
                   _d964, _d965, _d966, _d967, _d968}),
                    .FORW_LADDRAO({_d969, _d970, _d971, _d972, _d973, _d974, _d975, _d976, _d977, _d978, _d979, _d980, _d981, _d982,
                   _d983, _d984}),
                    .FORW_UADDRBO({_d985, _d986, _d987, _d988, _d989, _d990, _d991, _d992, _d993, _d994, _d995, _d996, _d997, _d998,
                   _d999, _d1000}),
                    .FORW_LADDRBO({_d1001, _d1002, _d1003, _d1004, _d1005, _d1006, _d1007, _d1008, _d1009, _d1010, _d1011, _d1012, _d1013,
                   _d1014, _d1015, _d1016}),
                    .FORW_UA0CLKO(_d1017), .FORW_UA0ENO(_d1018), .FORW_UA0WEO(_d1019), .FORW_LA0CLKO(_d1020), .FORW_LA0ENO(_d1021),
                    .FORW_LA0WEO(_d1022), .FORW_UA1CLKO(_d1023), .FORW_UA1ENO(_d1024), .FORW_UA1WEO(_d1025), .FORW_LA1CLKO(_d1026),
                    .FORW_LA1ENO(_d1027), .FORW_LA1WEO(_d1028), .FORW_UB0CLKO(_d1029), .FORW_UB0ENO(_d1030), .FORW_UB0WEO(_d1031), .FORW_LB0CLKO(_d1032),
                    .FORW_LB0ENO(_d1033), .FORW_LB0WEO(_d1034), .FORW_UB1CLKO(_d1035), .FORW_UB1ENO(_d1036), .FORW_UB1WEO(_d1037), .FORW_LB1CLKO(_d1038),
                    .FORW_LB1ENO(_d1039), .FORW_LB1WEO(_d1040), .CLOCKA({_d1041, _d1042, _d1043, _d1044}),
                    .CLOCKB({_d1045, _d1046, _d1047, _d1048}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na6948_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na6949_10, na6951_9, na6952_10, na6953_9, na6955_10, na6956_9, na6957_10, na6959_9, na6960_10, na6961_9,
                   na6963_10, na6964_9, na6965_10, na6967_9, na6968_10, na6969_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na6971_10, na6972_9, na6973_10, na6975_9, na6976_10,
                   na6977_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h000100906109030384018c330e9530023284c010240216c2300402184c208822000401084300f601),
             .INIT_01(320'h0753104000cf21c2c03d4c6100f531840004000000330870b00f61000100002012020081c2182080),
             .INIT_02(320'hcc2194649d6659d8660ce05040000080400242040f421b84300c1002000000324070a0c83a908219),
             .INIT_03(320'h8c3a1186208c6190040108c2181c318c188010000401081019874a580330e94308661d2f600cc3a5),
             .INIT_04(320'h8c61d0dc2104630e84e18823187433084118c3a1186208c61d0cc2104630e8461882318743308411),
             .INIT_05(320'h0c601ea62084019e43858660109630cf731806300f53184200cb6198c0318200400000803a138620),
             .INIT_06(320'hcc6018c03d4841000324870b0cc0212c61de8481cc6018c03d4c6100033c070a0cc0212c619ee630),
             .INIT_07(320'h0b1b04100000200ca33180630cc21c2c330084b186739843318063000324070a0cc0212c61de8481),
             .INIT_08(320'h807a98c201ea6308000800000cb21c0a0000401308421074100c617082208810104381e96200f430),
             .INIT_09(320'h0b520200800003ce839c2833c870b0e1780e043d084bc0f000e6781e8010003816200000019e4385),
             .INIT_0A(320'hef73d8943def63def4b1cf6310f4258c3a4cc421e841c8c7a167594005e57dc018f43d00228e8415),
             .INIT_0B(320'h0f41de061d0779c28321e801d014100401c0f021620040001004021080040f4bd0f63de84378c43d),
             .INIT_0C(320'h804200310000019eb601067a980419e96010661d041880000080401ef3a1bc001e039dc7385e7423),
             .INIT_0D(320'hebac00baaeb0031e85b5a9421884116a41cc520c4100400001873b0085a0e76010a41cec02128399),
             .INIT_0E(320'h8863dc873108620007b1886300e4210e4210f420e463d0bfafb8021715d600431e94a1a84148c7ae),
             .INIT_0F(320'h800004100004010040100402008c210b43108619084378843d29421287310943d2c7b909620007b1),
             .INIT_10(320'h07020013a408670ef330ef030ef330ef230ef130ef230ef130ef030e06610c03d284610c21c08c21),
             .INIT_11(320'h0709ce439982070607bd0de016501940385065210042708600e139c06599c749927719c761987419),
             .INIT_12(320'h62000000000403c3c190e6680e1419ec02908320871138303de84f00e380cd21c2c3290c021b8430),
             .INIT_13(320'h85c28421118c2e1846303863185c318c0e18c6130c613082301879182080002003c0082000006600),
             .INIT_14(320'h3848005c2401f80bc087612e821c84b8087a106124613092301849184c200c6130c4018c0e121231),
             .INIT_15(320'h80530b838184210bc1040001009090652002401480090a06198406104600820e1092070843000630),
             .INIT_16(320'h0020120c318208000201201170822008391000218c030842140431087010852010c214806300f02d),
             .INIT_17(320'h00420080210661d0c0218f5b100420ea7ad880210043d6c40108330ef530c83bd826014c02d82080),
             .INIT_18(320'h006618c1882000080330ef5b0cc021ec7ad8802100600cc3bd6c330087b1eb62008401803300f5b1),
             .INIT_19(320'h18421806300402185c2088220a04018208000201e86618c104000100003dcc0230c600e77394e6a1),
             .INIT_1A(320'h3a025ea597204bd2b0e009590002f045c248c0e100630bc28081e083d087820f400c318c2f085e84),
             .INIT_1B(320'h2000080400277a4806108301085c208822040410cb19c2b39d875850df87830f0097b165d812f5ac),
             .INIT_1C(320'h0c63004021204370c6300402138631842010dc318c010084e18c610804370c630040213c2618c608),
             .INIT_1D(320'h804210cc318c010084211863184201084330c63004021204230c63004021204370c6300402120437),
             .INIT_1E(320'h084b1867a8cc6018c330084b1867b98c031804214702800000cc0212c619666300c61c0a00004010),
             .INIT_1F(320'h0f23038381b863041000040078010400000cc00c4000000000800f0084203c0210840c4100000330),
             .INIT_20(320'h09230384018c0618803184c2424630185084223180c308c6170c6303863185c318c0e18c0e104617),
             .INIT_21(320'h2407824d001c0136007404e001b0032026000d009e0834127020d849d0838126c24c248c06124613),
             .INIT_22(320'h04411000200c330e8721b8630a41848329001200a429308230241130a480984210403185c24040e1),
             .INIT_23(320'h85290c121ca420480424812010c3346c10c41004000100933009c3180c3e1841104418080300c061),
             .INIT_24(320'h056300c221803b980421ab721480350c230886198c030cc0230c60044c20882200040c0843009204),
             .INIT_25(320'h09430843380c0e104411000206c335002018661d2b61d35481890310c3300c3b980421a972108035),
             .INIT_26(320'h840200c0100803d484010c010a420820000804830c60820000802008048025c2088220c040186601),
             .INIT_27(320'h8c03d0f7a1806300f4390c03184214cc021286008043980430840280c2900861009030840240c210),
             .INIT_28(320'h21437007b0467b0ee51de94850dc01ec11c0f02140080002012020c3841100408080210f43dc8601),
             .INIT_29(320'h0000000381e042820000800e805e003b017610e825e043b0082000007028000008033d87728ef4a5),
             .INIT_2A(320'h3b017800ec05d843b097813810f7010f421e9000e043dc043d20324073b0e821c0dd1c0dd1c0dd10),
             .INIT_2B(320'h3b097a06203b017610f40c417600ec25e81883a000081e803d240f02401c0b104000100e3a0270a0),
             .INIT_2C(320'h0403d09c318208000200007b9806e18c01cee729cd42009c31831040001005e80ec39c2c0f005d80),
             .INIT_2D(320'h802010d02138631802010dc318c210084e18c600804370c63084021386318020109e030c63041000),
             .INIT_2E(320'h084618c600804210cc318c2100842118631802010d021b8631802010d02138631802010d02138631),
             .INIT_2F(320'h0c33d464300c619804250c33dc86018c0210a381400000660109430cb32180630e05000020084021),
             .INIT_30(320'h070270c60820080002003c00820000066006200000000040078042101e0108420620800001980425),
             .INIT_31(320'h0803184c3100630184848c6130a10844630b86118c0e18c6170c6303863185c3185c208c0e1e4607),
             .INIT_32(320'h0401080010a02043840084c208c21044c2120261084100c61709010384901849184c248c06124617),
             .INIT_33(320'h040249863041000040281c4010041c880104100004010090a180021b86301c401004100801064210),
             .INIT_34(320'h8542168429086218443028600086618c0108800d4c00108c3184e2008220c4400e06104310401000),
             .INIT_35(320'h886110c3b9807cd90524006cdd0521c97210c430886110c21dcc0210d9ba0a4392e421886110c221),
             .INIT_36(320'h4e6a1006618c188200008020080499e6385c5e2008220e4409ec30005e2008220804010f31484430),
             .INIT_37(320'h0402138631842010dc318c010084f0b86318208000201e86618c104000100003dcc0230c600e7739),
             .INIT_38(320'h0848108c318c010084810cc318c010084810cc318c010084810cc318c010084618c610804330c630),
             .INIT_39(320'h0a00000330084a1865990c031870280001004201084330c63004021084618c610804210cc318c010),
             .INIT_3A(320'h62080002003c021080f0084210310400000cc02128619ea32180630cc02128619ee4300c6010851c),
             .INIT_3B(320'h0c061e06030860820000800f1004010222008698e701c0838104c21e80301843d080301843d08030),
             .INIT_3C(320'h2c2bd8402198430002f004c2c0c2610c20c410000403018430e6601086610c3998042198430e0661),
             .INIT_3D(320'h20314242010b01c001392e62139409085a1683a9094210049d604200949de04210020018430ec21c),
             .INIT_3E(320'h0901ca00988310400000802018061024050ef4010802027020e20e406284e4200084282000004210),
             .INIT_3F(320'h42588203948310401300000028020080210040feb0826ee461088441083d110421049de743c08421),
             .INIT_40(320'he95ab0879d10ce1384f14804611421aa7fd10420e610440210e000001c4111a02494250868008531),
             .INIT_41(320'h08427f2140318600845c0803de93a8eb440087a3f40c26c8e1086d708797084210442195c3d2c557),
             .INIT_42(320'h8021c088a1808e2b844a1f422042e30dc430f03200a21b839120421ac520ea3b6384370dc21084e1),
             .INIT_43(320'h0a021edc21384210862109fb10c0b70a003004211343d0a3ac40431087a108420000500401004010),
             .INIT_44(320'h18f4110c011042538437e84218842704437000e254022a40e0f001d05c000dc020942d0c421e8421),
             .INIT_45(320'h10950028624883d5b8c208810087a28960008b98042e1dc02228a2109c234dc418144118c7a10da1),
             .INIT_46(320'hef4010802027020e20612321000421410003f14111810b84418341eb8446040e6850630058b0eee1),
             .INIT_47(320'h44024000008002020000040100a427e0201177a0e041c44c90800210a08000010040100c02724042),
             .INIT_48(320'h09435ef53d884b5e941eee7a02e7bc49021a042108504010000400985021004240100000030bd01d),
             .INIT_49(320'h09041374ddf741e087a10f4a0cf6906100403421467c100000006013e480ee419ef7a70000080030),
             .INIT_4A(320'h04330880b9140bd2e7a02e781e93a04a5a40f41e0785dae33505799cda55b35c0025240902212544),
             .INIT_4B(320'ha7604ef714603c04f5000f480be835bd7a7882f92f6ea00705294a18f8e4b8459a9d50e801004010),
             .INIT_4C(320'h0004652824107be52881a0820ef421bf431bc401ac6f5876a000200802000c330a833d057d57783a),
             .INIT_4D(320'h403a06f8800f5803e4bd3f7a529c25ae411ad13d8f7b1e749cb9725e94e0b83b848621085a002812),
             .INIT_4E(320'h0f7ca510241041de9ea1b8435bc4118d6f98772000200802000c3308833d057d56f839a7a04ef714),
             .INIT_4F(320'h107a1000190193d2800c0421000811e960060040008028f4a00300287802102b20b6c1e83c950601),
             .INIT_50(320'h67441104b0084410082126288010220860c08784f8000b85a9917c6330ea0782229c07e81b8f7954),
             .INIT_51(320'h006000cc2212861084210843841094830000020d80200802000043000845ec04248801e882228610),
             .INIT_52(320'h8f4200eb2a4e40029d42167098082009d401794d106bdb884254c4108481086e00a8200004080210),
             .INIT_53(320'h0f7b68d631ed4b1b474a097c66d8a6ef4014e816cd739e54002a602080213a829f240017882f2441),
             .INIT_54(320'hef520863a0e87bc4f2010202009080004fa91c02005200173c48041806ea0f93d2e417f04c5f082d),
             .INIT_55(320'h20781000f92e4e508321c83a90001dea7008741d0f789e00240002001f25c9ca1064390752000205),
             .INIT_56(320'h05411a8019483b1e45b8af411e702d0179def024080fd480100763c88704a83c0077a024781017bd),
             .INIT_57(320'h002e0066bde44a82f4b9295b5ca4bdae5a5ed62508419a803d296392a0b1cc6b0494358e40d2e43d),
             .INIT_58(320'h085210862000011064803c6c6ec43ce96210a04100400004000942908417295a12802008010042e4),
             .INIT_59(320'h0803d4d42008620c8459074210041d2c400474310001d0441d0f4bd083b108021002fde943d0f420),
             .INIT_5A(320'h0b6a14802000390190200052c074208800128000804a0810110002106580c840100401004174801d),
             .INIT_5B(320'h1f4a1044130122001c720e7ae01fbd0843d4a827080008020080420233a00020c4100401c0008021),
             .INIT_5C(320'h0580108cc85b4e104c110401308420880250c419020250c419013a0087812f220c80138b001004b1),
             .INIT_5D(320'h728c2f6ad2728c2e62b16a4a1ee6b16a4a1e62b16a4a1ee6b16a4a1e629062080e62906208002c1d),
             .INIT_5E(320'h7ace3feef37ace3e62f37ace3feef37ace3e62d2728c2f6ad2728c2e62d2728c2f6ad2728c2e62d2),
             .INIT_5F(320'h5ad6ba800000000a800000000af7bdef7bdab5ad6b5adab5ad6b5ade62f37ace3feef37ace3e62f3),
             .INIT_60(320'he67514737807328df33bd7360ce379d8220c639906813a800000000a800000000a800000000aad6b),
             .INIT_61(320'hd211c46f79d811bd211c4233acf77acf33c46759de7dad011bd013dc6809ca3a9ce288e6f00d67ab),
             .INIT_62(320'hc0239ed300def3dce01102f98e641bd8339def38000000000000000000000033ddeb3cce379d811b),
             .INIT_63(320'hf46684781f077a046d6edeb3be8220de77ce812ec6414061b8e641a07a334201204c1946f60ca37b),
             .INIT_64(320'h12459cbf7d123db067329480420080a038dc7320d03d19a100031154310c8ce5245014e377cc8340),
             .INIT_65(320'hde6bdce01cdd3b9c663d46738053996fb990639d46f780040273b9c0500bcf334d833bce72800842),
             .INIT_66(320'heebd80773c46f99c012b64b1dcf6985e718e037cc6f195f734d6b1c066bd0663d00120e233847319),
             .INIT_67(320'h250b55697b461397fdde6f59c1cc520c410b9ec6a9684daf4aca7080473bd6d08df01402f1dd7b99),
             .INIT_68(320'h358f7461395697b6f59c7fdde0c4101cc52a9684b9ec6ca708daf4af3befe33ad90a6380221358f7),
             .INIT_69(320'h00000000000000000000000004bb99c4b008817df679906b3d06b3de33adf3bef8022190a63250b5),
             .INIT_6A(320'heefb9ee76caea7c0440bdf353d7320d0b99e6b39f63811990b680000000000000000000000000000),
             .INIT_6B(320'h1529cce5c0ac29cce5c09429cce5a0a4634e672d1575ce672d0671ac620d067bbeb01bea3acd8318),
             .INIT_6C(320'h080000001def73b1550fa2eb306748471808e7799301de7762dd35cce239c5819c6b9b60379ca2ac),
             .INIT_6D(320'h28798a418820398a41882000000000df41cd0379df01106339e6fbccec1bc6f68e651be0160e82c0),
             .INIT_6E(320'h30b98b49ca30bdab49ca30b98b49ca30bdab49ca30b98ac5a9287b9ac5a928798ac5a9287b9ac5a9),
             .INIT_6F(320'h6b798bcdeb38ffbbcdeb38f98bcdeb38ffbbcdeb38f98bcdeb38ffbbcdeb38f98b49ca30bdab49ca),
             .INIT_70(320'h002a000000002a000000002ab5ad6b5aea000000002a000000002bdef7bdef6ad6b5ad6b6ad6b5ad),
             .INIT_71(320'h023dc8c3749f048c733b075dbde788e23a8d8378ded1cca37c1777b0479dd7b9cc8340deea000000),
             .INIT_72(320'h000000733a023c9c8911c093bdbb51d601cd03d2c6c18e778088319cea38e641a1777b000000039a),
             .INIT_73(320'h0000000000003c8e691dcee1c02919f7790e0188c6e1c02f70e037c0780a4235cde942e755b003a0),
             .INIT_74(320'h00000000000000000000000000000000000000008000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6633 ( .DOA({_d1049, _d1050, _d1051, _d1052, _d1053, _d1054, _d1055, _d1056, _d1057, _d1058, _d1059, _d1060, _d1061, _d1062,
                   _d1063, _d1064, _d1065, _d1066, _d1067, _d1068, _d1069, _d1070, _d1071, _d1072, _d1073, _d1074, _d1075, _d1076, _d1077,
                   _d1078, _d1079, _d1080, _d1081, _d1082, _d1083, na6633_36, na6633_37, na6633_38, na6633_39, na6633_40}),
                    .DOAX({_d1084, _d1085, _d1086, _d1087, _d1088, _d1089, _d1090, _d1091, _d1092, _d1093, _d1094, _d1095, _d1096, _d1097,
                   _d1098, _d1099, _d1100, _d1101, _d1102, _d1103, _d1104, _d1105, _d1106, _d1107, _d1108, _d1109, _d1110, _d1111, _d1112,
                   _d1113, _d1114, _d1115, _d1116, _d1117, _d1118, _d1119, _d1120, _d1121, _d1122, _d1123}),
                    .DOB({_d1124, _d1125, _d1126, _d1127, _d1128, _d1129, _d1130, _d1131, _d1132, _d1133, _d1134, _d1135, _d1136, _d1137,
                   _d1138, _d1139, _d1140, _d1141, _d1142, _d1143, _d1144, _d1145, _d1146, _d1147, _d1148, _d1149, _d1150, _d1151, _d1152,
                   _d1153, _d1154, _d1155, _d1156, _d1157, _d1158, _d1159, _d1160, _d1161, _d1162, _d1163}),
                    .DOBX({_d1164, _d1165, _d1166, _d1167, _d1168, _d1169, _d1170, _d1171, _d1172, _d1173, _d1174, _d1175, _d1176, _d1177,
                   _d1178, _d1179, _d1180, _d1181, _d1182, _d1183, _d1184, _d1185, _d1186, _d1187, _d1188, _d1189, _d1190, _d1191, _d1192,
                   _d1193, _d1194, _d1195, _d1196, _d1197, _d1198, _d1199, _d1200, _d1201, _d1202, _d1203}),
                    .ECC1B_ERRA({_d1204, _d1205, _d1206, _d1207}),
                    .ECC1B_ERRB({_d1208, _d1209, _d1210, _d1211}),
                    .ECC2B_ERRA({_d1212, _d1213, _d1214, _d1215}),
                    .ECC2B_ERRB({_d1216, _d1217, _d1218, _d1219}),
                    .FORW_CAS_WRAO(_d1220), .FORW_CAS_WRBO(_d1221), .FORW_CAS_BMAO(_d1222), .FORW_CAS_BMBO(_d1223), .FORW_CAS_RDAO(_d1224),
                    .FORW_CAS_RDBO(_d1225), .FORW_UADDRAO({_d1226, _d1227, _d1228, _d1229, _d1230, _d1231, _d1232, _d1233, _d1234, _d1235,
                   _d1236, _d1237, _d1238, _d1239, _d1240, _d1241}),
                    .FORW_LADDRAO({_d1242, _d1243, _d1244, _d1245, _d1246, _d1247, _d1248, _d1249, _d1250, _d1251, _d1252, _d1253, _d1254,
                   _d1255, _d1256, _d1257}),
                    .FORW_UADDRBO({_d1258, _d1259, _d1260, _d1261, _d1262, _d1263, _d1264, _d1265, _d1266, _d1267, _d1268, _d1269, _d1270,
                   _d1271, _d1272, _d1273}),
                    .FORW_LADDRBO({_d1274, _d1275, _d1276, _d1277, _d1278, _d1279, _d1280, _d1281, _d1282, _d1283, _d1284, _d1285, _d1286,
                   _d1287, _d1288, _d1289}),
                    .FORW_UA0CLKO(_d1290), .FORW_UA0ENO(_d1291), .FORW_UA0WEO(_d1292), .FORW_LA0CLKO(_d1293), .FORW_LA0ENO(_d1294),
                    .FORW_LA0WEO(_d1295), .FORW_UA1CLKO(_d1296), .FORW_UA1ENO(_d1297), .FORW_UA1WEO(_d1298), .FORW_LA1CLKO(_d1299),
                    .FORW_LA1ENO(_d1300), .FORW_LA1WEO(_d1301), .FORW_UB0CLKO(_d1302), .FORW_UB0ENO(_d1303), .FORW_UB0WEO(_d1304), .FORW_LB0CLKO(_d1305),
                    .FORW_LB0ENO(_d1306), .FORW_LB0WEO(_d1307), .FORW_UB1CLKO(_d1308), .FORW_UB1ENO(_d1309), .FORW_UB1WEO(_d1310), .FORW_LB1CLKO(_d1311),
                    .FORW_LB1ENO(_d1312), .FORW_LB1WEO(_d1313), .CLOCKA({_d1314, _d1315, _d1316, _d1317}),
                    .CLOCKB({_d1318, _d1319, _d1320, _d1321}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na6985_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na6986_10, na6987_9, na6989_10, na6991_9, na6993_10, na6994_9, na7000_10, na7002_9, na7005_10, na7012_9,
                   na7013_10, na7016_9, na7030_10, na7035_9, na7037_10, na7045_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7048_10, na7050_9, na7053_10, na7056_9, na7058_10,
                   na7060_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h018a5002e020021982c300621f822150020886a1f0400885c1284080fb20a0020cd8000022104020),
             .INIT_01(320'h0040818520a8c6100c010006100404185000f0040032018403804612003c01060030240d0120841c),
             .INIT_02(320'h805c500411024110440108020e0083180010102007c20102418042107004002a1184030802050c21),
             .INIT_03(320'h004204000148021082400641208809004210838020c04080110fc1109221f82213c43f0402b887e0),
             .INIT_04(320'h88021030040bc0108220185a00840d00c29004207004148021010020a40108360085200841100429),
             .INIT_05(320'h10421080850b091194a02c422102010fc300882108400285840c42180441084a4c00831802040081),
             .INIT_06(320'h0c022084010288171221214048844204021f83e00c022084210208171223294058844204021f8601),
             .INIT_07(320'h002210934041ce00843008821a806100e211081008601184300882158221214048844204021f81e0),
             .INIT_08(320'h1802020c20080030a001e004088421007c03141c00042b06c31803dc8280d815a00c200816007c0c),
             .INIT_09(320'h067262949a0100368c0100ea0104020806208c6018c0320d20084600847000020087802001518c20),
             .INIT_0A(320'hfe821e037fd67bfd741d087bc00760e9ba00f01be800100020004030000200c00efc1a30020d0019),
             .INIT_0B(320'h0043f008391fc0100c2008461080660480100400084a4d00c4297400002007c010079fd0002df01f),
             .INIT_0C(320'h180010043c00801f8003087e000821f80010841f08421f00c528008f87e0a042001be100c2018408),
             .INIT_0D(320'h000600006018019f8339082afa8015ad5865294a52528a00801842318001084620002108c2000421),
             .INIT_0E(320'hc82810e03903ea008034c8290c06e0a8700ad4000800100020180000080300015f8015c800100020),
             .INIT_0F(320'h080040930061d084a54a5ae80064180645506021c0016adc1f002a4055b9002b906421b832008034),
             .INIT_10(320'hf148008020001c1295c1295c1495a1495c1695c1695a1895a1895a1283e01041f000e0104e501c02),
             .INIT_11(320'h394012f4ad08f61003e30582000079014a02f4062801a00827280257d4c1045a56c64595739cd7c9),
             .INIT_12(320'h087c00000041c05e04022e4042808d087a0313e4314070801f1806100003c8085013a03100030041),
             .INIT_13(320'h0dc0000009004a002401902200d00f006e0680200083b00041b83e20849801060c84010700200421),
             .INIT_14(320'ha80002a4002b800780110024005000a8017000600002b00001a000008c161803206003004e000120),
             .INIT_15(320'h0808128020b04a148024d0107001c123c20885520ae8141025006a000033085a0800540000228421),
             .INIT_16(320'h01060068020841c018a0004117012048103000002041d0d42cb85b80b74166c200182908081a0c04),
             .INIT_17(320'h00180000820143f02c000041f0018008020f800c0000107c00600a1ffc81683e101034205840841c),
             .INIT_18(320'h082201042126804180a1ffc812844208020f800c0102b287ff204a110820083e0030040d8a10041f),
             .INIT_19(320'h6800408c01904040b9c04822073c040849a01060f802010420e00c50039f08c0a008200840100400),
             .INIT_1A(320'hf8000f80620001f00cc000078000c10800000780b0c01684130c021a80130ff0004809007012f400),
             .INIT_1B(320'h0700628001007e01806a091811c9c0482209cc032886100c21184600281308300003e01ec0007c03),
             .INIT_1C(320'h0240128400a000302401b0400001200e82005809007e1001a0480230800302401e84004068048021),
             .INIT_1D(320'h08042014110066100840581e00e0201081003401984001000102401c84004001f02401f840070001),
             .INIT_1E(320'h10804087e109022084a110804087e1204410884108401f004028442010210848110421007c020c0d),
             .INIT_1F(320'h07c41b00a0a00410930020c1908020e0040084210f800000041806100841304021082108380100a1),
             .INIT_20(320'h00001782c3007c0c00600c8000240118000001200c4004803d04401001e00880d00580104e000822),
             .INIT_21(320'h010000040018404080c001c0048015002c006020c801b0038107820f80010004003800006e00003f),
             .INIT_22(320'h0140402460204a10c3c0c0041704900822154c2ba051100001f042900c0280000110210c400010c0),
             .INIT_23(320'h0b0a169c2d4058a080020e020006a0f0422314a4d0107000a10140208c00024050100950381e04e9),
             .INIT_24(320'h004a1304e70b0a5080000882010001304a139c29284c1284040083f0792028220730000000106424),
             .INIT_25(320'h103c1a85b1f05a90141104640f04a50003c0f43f0782de340008007384a1304a5080000842008001),
             .INIT_26(320'h70400f052100c0105c00f066102c2107004180070082107006190852800100120282208e01e0f422),
             .INIT_27(320'h0841f007e00882107c01004410d020e84420783408181083c110400f04c100241007c150400f0541),
             .INIT_28(320'h08015030210b421f843f080200780c08421004000841c0106006424f240500016d800007c01f8022),
             .INIT_29(320'h2100021020080012600418100024205800c001c003c20884010700200401f0083181a10fc21f8400),
             .INIT_2A(320'hf84000804000c0028406080a2104a217c42080a72884128841014a01842309081038250402504821),
             .INIT_2B(320'hf80000018018004000c0030080014002c00601a0004000840100e8006c0100424d0107017a509405),
             .INIT_2C(320'h20c1f04c020841c018a0073e11836010401080200800100c0208424d00c505c0028c0100f8007400),
             .INIT_2D(320'h0942004800101200d8200780900741002a04803f0800b0240118400101200f420054330240108380),
             .INIT_2E(320'h1008088033080420240f0070100840781a00cc2000000f81200e42001800f01200fc200300000120),
             .INIT_2F(320'h0043f0840110421088400043f0802208442084200f802004221000108420088210803e0106068402),
             .INIT_30(320'h01412008212949801060c84010700200421087c00000020c030804209820108410841c0080108840),
             .INIT_31(320'h058600ec1800c018000048020000000240170009007608803d03c01001a00a4020900010400f8835),
             .INIT_32(320'ha05550aee147820d8000220000048108010008e0000440842800004e8004600000d000007a00002c),
             .INIT_33(320'h20c00c80410838020c0082c0703c07601c108380418e7000a5080003004102c07018062022124820),
             .INIT_34(320'h1b40008011000e71a1034a4600036010fc32000630c0000c021f160382204bc0528283099494a2c0),
             .INIT_35(320'h4206738d29180210802000021080200080011ce34206a50e0948c000042100400100024206738d4a),
             .INIT_36(320'h0040008260104212680a3a10948015f94a02d960382205dc0b08ca927960382205cc00004210a943),
             .INIT_37(320'hf8400e012008c2004809007a1002a1181200841c01060f806010420e00c50039f08c0c0082008401),
             .INIT_38(320'h002200400900721002e003809007e1003a004009004a10006004809006c1001e04803a0800502401),
             .INIT_39(320'h007c0101211080b084215844108401f00830342010814044019840210340780380804207c0d00661),
             .INIT_3A(320'h0849a0106018402104c10084208420e00404844202c21f842b088214844202c21f85611042210421),
             .INIT_3B(320'h205409902701021268062822b01c1c04f200006318421084220f400f84810801f084812801f10481),
             .INIT_3C(320'h00d211840008081380a10c401205c0204210934031403e808108460102802042118020c808108380),
             .INIT_3D(320'h318a5010af01405c002100442e800100020083e1e00000701f08000e001f00000018a038081c8061),
             .INIT_3E(320'h00c6211482108c5d0144214a010061080070fc0100000086c00800a524a44806000006296c040ee1),
             .INIT_3F(320'h080eb5ad4a529cd6b152018800042210c64296b6174c0f8820000140001f060000002307c0400000),
             .INIT_40(320'h08060020bfd4762e07a006700000000813fe2782794a16b5cd18000068140000300060c008007000),
             .INIT_41(320'h00212cbf2118c2000440083e08b020fcc8010ae0aa6d2745288206b0142d00080e00083c88100815),
             .INIT_42(320'h635bfe0000007a000022efc80200800780007d000000058c20000000900008bf38001184800002b0),
             .INIT_43(320'h80442ee442d8c6007000050600202500468001001045d004210802007c0c0420073007421295296b),
             .INIT_44(320'h10be8420081205dd085bf801c000100000d006e00018020262a89617d9e21306217e810801f04014),
             .INIT_45(320'h00000988011300d10c04200c040021d002160021202d801800084400018107000100081085d00060),
             .INIT_46(320'h0fc0100000086c0082402180300000314b8bf44c00080830000087fa40003032001400200a0a03b8),
             .INIT_47(320'h0cc000f8020ab9507806210a50040408400007e00d8010748018000018a5d0105318e70081608000),
             .INIT_48(320'h083011fc43084011801f08424025a30a8005801005041083c0100210e80028001083c010401d8401),
             .INIT_49(320'hff8000fc3f17c2200020d7cdfffc4210420f8400107e0e00020842118401087c108c7c0004000401),
             .INIT_4A(320'h18c202881108022080000842108065087eb0650d007010842127465088410800040420fe80000420),
             .INIT_4B(320'hffc4008842107e10fc400083c485095d62d781df04601f97e008000004c0b81416e8200808008442),
             .INIT_4C(320'h00420087e1003e20841f28000f8a1098781abc140870200440200010884300c202fc3f017e10fc01),
             .INIT_4D(320'h317e10fca00085adfc1dd84410c80028401084210847918409d0030182c05fcbf810400044c00401),
             .INIT_4E(320'h07c41083e10001f148209f015abc1508702004403084319085014202fc3f077e10fc01ffc4408842),
             .INIT_4F(320'h180a01441f0002305401006e100001183600801e0000010c020040020400000420984a087e10ff80),
             .INIT_50(320'h08403108670000250800198c629000000c618c45f8078e84411004108b21e0800078070fcdf7fc23),
             .INIT_51(320'h1806003c00005400218000002104021083c020c110c64214a638007d000117002083e20806218823),
             .INIT_52(320'h0fd14084210848003441604613800902c3d004210103f780000e40001000a02e0004002080000422),
             .INIT_53(320'h00fe1088221840108441080600840018c000840108435184042064005000b84210848b0640008408),
             .INIT_54(320'h088210cc210fca208c800040000021f51e208480001a0201230c80098121084210051a084001c201),
             .INIT_55(320'h003e0002bf056e00802308421080411066108421f94411c0000fa00053e0ad801004610842100801),
             .INIT_56(320'h004400800168021104220fc25f8d09043ff17c00003a168041c0422288400fbe107d200046c043e2),
             .INIT_57(320'h0f260004210840007c01000010800108400f84001080108001000210000108420003c10842000401),
             .INIT_58(320'h00025034000000500400d0c6229801780d8001a00040001800600001081c00020000000008108e20),
             .INIT_59(320'h28305885a0200000971fc74a80040f01400084c6000190180503c01683a6200c100325780a1804a0),
             .INIT_5A(320'h0842d0000000be10007e000a0074a028018060020e01840008f00960040008804010040101c08015),
             .INIT_5B(320'hd040e0001d0817e06c24c07e1c583f000010141f0008108843191a000020c604210420e4c0000000),
             .INIT_5C(320'h0100739ce739d0a0005b0042310ac0103800040100380004010002010ba007000080158800906000),
             .INIT_5D(320'h08421000000000008421084210000000000084210842100000000000842108421000000000000803),
             .INIT_5E(320'h08421000000000008421084210000000000084210842100000000000842108421000000000008421),
             .INIT_5F(320'h00000100000000010842108421042108421100000000010421084210842108421000000000008421),
             .INIT_60(320'h01018449c40425252812400c046246f03c0048ca0701810000000001000000000108421084210000),
             .INIT_61(320'h0394a10b400014e0394a1100804148c191060100a029c4014a4010a3200846248320489388007200),
             .INIT_62(320'h20100428801680c0201e0188a3281a70100d380400000000000000000000000105230646b400014e),
             .INIT_63(320'h5100c123ca009805280052808d03c072b0af02004001c0000632808028806081802812309409184e),
             .INIT_64(320'h0234a00108a481eefbe4315c11bc40e0004319404014403058043ca94250411064081c0700650100),
             .INIT_65(320'h9008a02002229404009e378080201c410ca01900409c4038c002a9a07006c1940103044308805152),
             .INIT_66(320'h068040021c42940202008238a7190600246403ca508c0060ca570c80508a0508a0020052bc044808),
             .INIT_67(320'ha52b594a73842317bdce6b58c5ad4a4a50839cc62948418c420840007812400905281c019dad00ca),
             .INIT_68(320'hbded68c6109ce52631ad739ef421295296b210a5318e70002110863f7bffe73bdd6b7bc6339b5af7),
             .INIT_69(320'h00000000000000000000000008014a320c0f00ca368ca02b4a02b4aef79cfffdece718def5aad694),
             .INIT_6A(320'h46a4000114109230780652a02319404010007b84520c739ce7380000000000000000000000000000),
             .INIT_6B(320'h0110051a80a210051a80a210051a80848c8028d40098af28d4050c68609405140050080205400100),
             .INIT_6C(320'h3800000002603480694a4034a020d2710c0a19c2e1000d73c0f0b92c180685014173c010140c4040),
             .INIT_6D(320'h000210842108400000000000000000508085010ac201e00384501865000ad29408494a5004018080),
             .INIT_6E(320'h00021084210840000000000210842108400000000002108421084000000000021084210840000000),
             .INIT_6F(320'h08421084210840000000000210842108400000000002108421084000000000021084210840000000),
             .INIT_70(320'h00040000000004210842108400000000040000000004210842108410842108440000000004108421),
             .INIT_71(320'h02814c010a3280a3201c05004001065011a0015a528109294a00b000781cd0186501005284000000),
             .INIT_72(320'h00000019080501020142303185035cd1008500083000640080f001c22b0a3280800b00000000010a),
             .INIT_73(320'h00000000000028a018925734a05200a281a5028a45b4a0725a501520281454bc051a800001e00300),
             .INIT_74(320'h0000000000000000000000000000000000000000f800000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6634 ( .DOA({_d1322, _d1323, _d1324, _d1325, _d1326, _d1327, _d1328, _d1329, _d1330, _d1331, _d1332, _d1333, _d1334, _d1335,
                   _d1336, _d1337, _d1338, _d1339, _d1340, _d1341, _d1342, _d1343, _d1344, _d1345, _d1346, _d1347, _d1348, _d1349, _d1350,
                   _d1351, _d1352, _d1353, _d1354, _d1355, _d1356, na6634_36, na6634_37, na6634_38, na6634_39, na6634_40}),
                    .DOAX({_d1357, _d1358, _d1359, _d1360, _d1361, _d1362, _d1363, _d1364, _d1365, _d1366, _d1367, _d1368, _d1369, _d1370,
                   _d1371, _d1372, _d1373, _d1374, _d1375, _d1376, _d1377, _d1378, _d1379, _d1380, _d1381, _d1382, _d1383, _d1384, _d1385,
                   _d1386, _d1387, _d1388, _d1389, _d1390, _d1391, _d1392, _d1393, _d1394, _d1395, _d1396}),
                    .DOB({_d1397, _d1398, _d1399, _d1400, _d1401, _d1402, _d1403, _d1404, _d1405, _d1406, _d1407, _d1408, _d1409, _d1410,
                   _d1411, _d1412, _d1413, _d1414, _d1415, _d1416, _d1417, _d1418, _d1419, _d1420, _d1421, _d1422, _d1423, _d1424, _d1425,
                   _d1426, _d1427, _d1428, _d1429, _d1430, _d1431, _d1432, _d1433, _d1434, _d1435, _d1436}),
                    .DOBX({_d1437, _d1438, _d1439, _d1440, _d1441, _d1442, _d1443, _d1444, _d1445, _d1446, _d1447, _d1448, _d1449, _d1450,
                   _d1451, _d1452, _d1453, _d1454, _d1455, _d1456, _d1457, _d1458, _d1459, _d1460, _d1461, _d1462, _d1463, _d1464, _d1465,
                   _d1466, _d1467, _d1468, _d1469, _d1470, _d1471, _d1472, _d1473, _d1474, _d1475, _d1476}),
                    .ECC1B_ERRA({_d1477, _d1478, _d1479, _d1480}),
                    .ECC1B_ERRB({_d1481, _d1482, _d1483, _d1484}),
                    .ECC2B_ERRA({_d1485, _d1486, _d1487, _d1488}),
                    .ECC2B_ERRB({_d1489, _d1490, _d1491, _d1492}),
                    .FORW_CAS_WRAO(_d1493), .FORW_CAS_WRBO(_d1494), .FORW_CAS_BMAO(_d1495), .FORW_CAS_BMBO(_d1496), .FORW_CAS_RDAO(_d1497),
                    .FORW_CAS_RDBO(_d1498), .FORW_UADDRAO({_d1499, _d1500, _d1501, _d1502, _d1503, _d1504, _d1505, _d1506, _d1507, _d1508,
                   _d1509, _d1510, _d1511, _d1512, _d1513, _d1514}),
                    .FORW_LADDRAO({_d1515, _d1516, _d1517, _d1518, _d1519, _d1520, _d1521, _d1522, _d1523, _d1524, _d1525, _d1526, _d1527,
                   _d1528, _d1529, _d1530}),
                    .FORW_UADDRBO({_d1531, _d1532, _d1533, _d1534, _d1535, _d1536, _d1537, _d1538, _d1539, _d1540, _d1541, _d1542, _d1543,
                   _d1544, _d1545, _d1546}),
                    .FORW_LADDRBO({_d1547, _d1548, _d1549, _d1550, _d1551, _d1552, _d1553, _d1554, _d1555, _d1556, _d1557, _d1558, _d1559,
                   _d1560, _d1561, _d1562}),
                    .FORW_UA0CLKO(_d1563), .FORW_UA0ENO(_d1564), .FORW_UA0WEO(_d1565), .FORW_LA0CLKO(_d1566), .FORW_LA0ENO(_d1567),
                    .FORW_LA0WEO(_d1568), .FORW_UA1CLKO(_d1569), .FORW_UA1ENO(_d1570), .FORW_UA1WEO(_d1571), .FORW_LA1CLKO(_d1572),
                    .FORW_LA1ENO(_d1573), .FORW_LA1WEO(_d1574), .FORW_UB0CLKO(_d1575), .FORW_UB0ENO(_d1576), .FORW_UB0WEO(_d1577), .FORW_LB0CLKO(_d1578),
                    .FORW_LB0ENO(_d1579), .FORW_LB0WEO(_d1580), .FORW_UB1CLKO(_d1581), .FORW_UB1ENO(_d1582), .FORW_UB1WEO(_d1583), .FORW_LB1CLKO(_d1584),
                    .FORW_LB1ENO(_d1585), .FORW_LB1WEO(_d1586), .CLOCKA({_d1587, _d1588, _d1589, _d1590}),
                    .CLOCKB({_d1591, _d1592, _d1593, _d1594}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7069_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7070_10, na7073_9, na7074_10, na7075_9, na7077_10, na7079_9, na7080_10, na7081_9, na7083_10, na7084_9,
                   na7085_10, na7087_9, na7088_10, na7089_9, na7091_10, na7092_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7093_10, na7095_9, na7099_10, na7101_9, na7103_10,
                   na7104_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h00000001603000048080000200002000000080802000008020180010314050160030000002000400),
             .INIT_01(320'h0000000000780000000000000000000000003c00001e000000080000000f0000000000024010000f),
             .INIT_02(320'h080000000000000000000000078000000000000000000480200800003c00001e0000000000000000),
             .INIT_03(320'h0000040000000000002003c010340000000001e00000500001000010002000020004000040008000),
             .INIT_04(320'h00000020000000000100000000000e00000000006800000000030000000000140000000000900000),
             .INIT_05(320'h00000000000000f00000004000002000001000000000000000004000800000000780000000040000),
             .INIT_06(320'h004000000000000001e0000000800000400000e0004000000000000001e000000080000040000020),
             .INIT_07(320'h00020001e0000000000100000780000002000001000200000100000001e0000000800000400000e0),
             .INIT_08(320'h000000000000000000007800008000001e00000900000200800000c501406002c000000014000000),
             .INIT_09(320'h03de00000f0000078000001e00000000000010002000000000000000000000000001e00000f00000),
             .INIT_0A(320'h7bc00781ef7bdef7bc0f001ef001e0781e003c0f78004000000000000000000007bc0f080007800f),
             .INIT_0B(320'h0000f0000f03c0000000000000000000000000000000078000001e00000000004001ef7800e7bc00),
             .INIT_0C(320'h000000000f00000000000000000000000000000000000780000000f001e06800000000000000000d),
             .INIT_0D(320'h00000000000000f781ef001e17800f7bc00000000000078000000000000000000000000000000000),
             .INIT_0E(320'h781e003c0f005e00000f781e0781e0781e07bc00200000000000000000000000f7800f7800400000),
             .INIT_0F(320'h00000001e00000000000001e00200f03c0f03c00780097bc00001e003def001ef03c00781e00000f),
             .INIT_10(320'h001e0000000012000020000200002000020000200002000020000200010000000001400000002400),
             .INIT_11(320'h00000000010010000000024000000f0000003c000000f00000000000800000400004000040000400),
             .INIT_12(320'h001e000000000007800003c0000001001e0001e00000800000001200000078000001e00000078000),
             .INIT_13(320'h0340000000001a0000004800002400001200000f0000f00000781e00000f00000781e003c0000000),
             .INIT_14(320'h5800002c0003c007800f001e003c007800f00120000090000048000038040000c02400001e000000),
             .INIT_15(320'h000006800018020680007800000000000000000000000000000010000003001e07800e0000000000),
             .INIT_16(320'h0000002c000000f000000000e681a06800d000000000201c0038007000e00000000c000000000000),
             .INIT_17(320'h000010040008000004000000c00001200006000008000030000040003c000040400001000200000f),
             .INIT_18(320'h001400000003c000000003c00000002000060000080000000f00000000800018000020000000000c),
             .INIT_19(320'h40000000002000002da0681a0034000000f00000781400000078000001e00000a000000100001000),
             .INIT_1A(320'h480000000a000000014000000001c002c00001e02000070001038005000e0014003800001c00a800),
             .INIT_1B(320'h03c0000000001e00000200060025a0681a0034007800000000000000240d00120000000240000000),
             .INIT_1C(320'h00000100000800d0000008000680000040002c000002000140000020000900000100006818000000),
             .INIT_1D(320'h0000002400000000000048000000000000900000080000800900000080000800e00000080000800e),
             .INIT_1E(320'h0000000000000000000000000000000000000000000007800000000000000000000000001e000000),
             .INIT_1F(320'h03c007800058000001e00000f03c00780000000003c0000000001e0000007800000000001e000000),
             .INIT_20(320'h0000048080001e04800002800000004800000000020000000c00000680000340000140001600000b),
             .INIT_21(320'h0016002c005800b0016002c005800a00140028005000a00140028005000b0016003000001800000c),
             .INIT_22(320'h004010002000000025e0400002000400080010002000b000000800a01800480000000003800001c0),
             .INIT_23(320'h0006000c00180040000100c001000008000000007800000000020000244050401004000802008141),
             .INIT_24(320'h0100000000000000000000000000040000000000000000000f000010202008020004000004000003),
             .INIT_25(320'h0002000000081e100401000200800000001004000040008000000000000000000000000000000000),
             .INIT_26(320'h08000080800000003400080a00180003c000000c0000003c00000000000003c20080200040100400),
             .INIT_27(320'h00000001e20000000000100000100008000004070002000020080000800000040000200800008040),
             .INIT_28(320'h0000b0040000400000000000002c0100000000000000f00000018006040100800080000000078800),
             .INIT_29(320'h00000000000000003c000016002c005800b0016002c005800003c000000078000000200000000000),
             .INIT_2A(320'h4800a00140028005000a000040000403c80000000100001000000000000000000028000280002801),
             .INIT_2B(320'h4000900001480090012000029001200240000401000000000000120000000000078000001c000000),
             .INIT_2C(320'h0000f038000000f0000003c00001c000000200002000003c00000007800002000780000010002000),
             .INIT_2D(320'h0080000000600000040002c00000200014000001000090000010000400000080003c0b00000001e0),
             .INIT_2E(320'h00100000000000002000000000000040000004000000078000004000000068000004000000068000),
             .INIT_2F(320'h100000004000002000001000000800000000000003c00008000004000002000000000f0000000000),
             .INIT_30(320'h0000a000000000f00000781e003c0000000001e0000000000f0000003c00000000000f0000200000),
             .INIT_31(320'h0100003809000004800000008000000000078000001600000b00000600000240002800001407800f),
             .INIT_32(320'h30006000c000c006800002c00000800280f00120000000000e00000680005800002c000016000008),
             .INIT_33(320'h0000070000001e000000488020080010000001e0000000000000000400005080200800100c001800),
             .INIT_34(320'h0000000000000000000000000001c0000e0180000000003c00020401004000800000e000000001e0),
             .INIT_35(320'h00000000000000000000000000000021000200000000000000000000000000004200040000000000),
             .INIT_36(320'h01000001800000003c00000000000f18000038401004000800000000384010040008000000000000),
             .INIT_37(320'h0800070000008000340000040001e0480000000f00000781800000078000001e00000c0000001000),
             .INIT_38(320'h000a00340000020000a002c0000020000a00280000040000c0024000002000120000010000800000),
             .INIT_39(320'h001e0000000000000000000000000078000000000000d0000000000001a000000000000340000020),
             .INIT_3A(320'h0000f0000078000001e0000000000078000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h001c00000d0000003c00001220080200040000000000000000038000000078000000007800000000),
             .INIT_3C(320'h000000000068000001c0034000018000000001e0000006000000000001a0000000000068000001a0),
             .INIT_3D(320'h00000000040000078000000007800400000001e47800003c0f000007800f00000000006000078000),
             .INIT_3E(320'h1000000000000007800000000000200000003d0002000001a0001e0000000000000000001e000020),
             .INIT_3F(320'h0000000000000000000f000000000000000001ef03c0000000000000000000000000040340000000),
             .INIT_40(320'h0000000000781e0781e0001e000000000007806000000000000000003c0200000000001000000800),
             .INIT_41(320'h1000f701c42002008060001e00000003c00001e000000001e00800f0008f000000000003c000000f),
             .INIT_42(320'h0000f70000001e0780807bc00001e00280003c03000007800000000010001000f7000e13822005c0),
             .INIT_43(320'h000007bc807900013c000bc800048b00001000000000f210840000003c0010000000000000000000),
             .INIT_44(320'h001e003c0f0000f7800f0004f0002f0000f00160001c0001e07880003c0003c0003c000000f00040),
             .INIT_45(320'h0000000004000002000068000000047800068000001ef20000010000000003c00000000000f00000),
             .INIT_46(320'h03d0002000001a0001c000000000000000f4bc8c0000063c000000f63c00001e000004000007918f),
             .INIT_47(320'h0040003c00005e103c00000000000800000001e80340003400000000000078000000000000800000),
             .INIT_48(320'h001e403c04200000000f0008000000218003000000000001e00000401c0000000001e00000078000),
             .INIT_49(320'h790000000003c00000000bc277bc000000038000001e07a0000100078000211e00108f0000000000),
             .INIT_4A(320'h000000000000000000000000400000201e4000000100000004000002000000008010007900001000),
             .INIT_4B(320'h03c0000000001e0000080000f781ef7bdef201ef03de03bc0000000001e07800003c000000000000),
             .INIT_4C(320'h40000011e2000002000f10000001ef781e07900f001e00000000000000000000001c0f405e000000),
             .INIT_4D(320'h001e0000080000f7bc0f780000380000100000000000e010007800f001e079c00780000000300000),
             .INIT_4E(320'h00004001e00000003c007bc0f7900f001e00000000000000000000001c0f405e00000003c0000000),
             .INIT_4F(320'h000000000f000000000400000000000000020000000000000101000080000008000c87001e003ce0),
             .INIT_50(320'h00000000070000038000000000000000000000007800f6800000000039e4380000380e01c0003c80),
             .INIT_51(320'h0000003800001c00000000000000000000f000000000000000000003000001800000c00000000007),
             .INIT_52(320'h03c20000000100003c00780042000403c04000000000f780000340000000001e0000000000000000),
             .INIT_53(320'h001e40008021004000840000000000000000000000080004000106000c0070000010040380000000),
             .INIT_54(320'h000800000003c00200404100000000781e003c00001c0001c020800101e0000000100d00000001e4),
             .INIT_55(320'h001e0001ef03de00200000004000000100000000780040040003c0003de07bc00400000008000000),
             .INIT_56(320'h0100000000780040000003c007800003de003c00001e078000080800000003de003c080000003c00),
             .INIT_57(320'h03d20000002100003c000000000000000000000000000000040000400000000800000001000001e0),
             .INIT_58(320'h0000040101785e00a00f78000000000000f000080a02f7802000000421ef00000000000000000120),
             .INIT_59(320'h00160000010010f0016f5bc000806000020010000840f0000000000005e00040008de00000000000),
             .INIT_5A(320'h0000100463001e05806f0000003c010040b02c0002c0b000087800a0200f421e0080200802f43c0f),
             .INIT_5B(320'h48003021e90006f03d43581e05bc0f000000000b000000000000020000015bc00000007bc0018060),
             .INIT_5C(320'h0000000000001e302403000090006043de0021e8789e0021e87890f001e003d0f40de91800300008),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h11c46398c7018c631806388e0318c730080398c60180400000000000000000000000000000000000),
             .INIT_61(320'h11c46318c23804611c4631447018c711cc6208e01806638046380c631c06398c6398c7318e0118c2),
             .INIT_62(320'h38062398e03184611804018e6318063006231847000000000000000000000000631c47318c238046),
             .INIT_63(320'h1144421064018a011c4231c4710080318c7200a23880401c6631807008a22100401006298c0314c6),
             .INIT_64(320'h39866108c70004520c642108421080200e3318c0380451108301c8421c872148420c04008e6300e0),
             .INIT_65(320'h300e611806398c2300e6298460140218cc601ce0298c7000001086501006318c0300c7318e700040),
             .INIT_66(320'h018e7008e6318c2380a2390c631ce7108c7380c6318e2118e7318e700ce600ce6000a0310c0218e6),
             .INIT_67(320'h100c45a5ed184e56390a218026bd2b29c2373148310407b5693946101006388c631804018c631cc6),
             .INIT_68(320'h5a5ed100c4521cc29c236bd2b218026390a394617b56931040731484298e008864adaf08ca7521cc),
             .INIT_69(320'h7bdef781ef7bdef7bdef7bde0388c6390e0200c6318c6018c7018c708ca74adaf008864298e184e5),
             .INIT_6A(320'h218c2108e30000001006318e6398c0380e2118c721cc000000001ef7bdef7bdef7bde07bdef7bdef),
             .INIT_6B(320'h014a231c60014a231c60014a231c60210a5118e3010e6318e3000e7318a3000c210c07114c3000c2),
             .INIT_6C(320'h00000000062806700ca228864018c639c6001cc630c00198a0310c61184738c00318c2180c231883),
             .INIT_6D(320'h00000000000000000000000000000039807300c631c0401cc7214a63000731cc2318463000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00843308e629c0239c4600046108e531ce6000e639846308c6018c20100231cc6300e03980000000),
             .INIT_72(320'h0000001cc70004738044380c6388c631c073004438007388e0200e6390c631807018c200000000e6),
             .INIT_73(320'h00000000000000211ca63988600042198443000239886008c4300c601802118c731c4010806000c0),
             .INIT_74(320'h00000000000000000000000000000000000000003842100000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6635 ( .DOA({_d1595, _d1596, _d1597, _d1598, _d1599, _d1600, _d1601, _d1602, _d1603, _d1604, _d1605, _d1606, _d1607, _d1608,
                   _d1609, _d1610, _d1611, _d1612, _d1613, _d1614, _d1615, _d1616, _d1617, _d1618, _d1619, _d1620, _d1621, _d1622, _d1623,
                   _d1624, _d1625, _d1626, _d1627, _d1628, _d1629, _d1630, na6635_37, na6635_38, na6635_39, na6635_40}),
                    .DOAX({_d1631, _d1632, _d1633, _d1634, _d1635, _d1636, _d1637, _d1638, _d1639, _d1640, _d1641, _d1642, _d1643, _d1644,
                   _d1645, _d1646, _d1647, _d1648, _d1649, _d1650, _d1651, _d1652, _d1653, _d1654, _d1655, _d1656, _d1657, _d1658, _d1659,
                   _d1660, _d1661, _d1662, _d1663, _d1664, _d1665, _d1666, _d1667, _d1668, _d1669, _d1670}),
                    .DOB({_d1671, _d1672, _d1673, _d1674, _d1675, _d1676, _d1677, _d1678, _d1679, _d1680, _d1681, _d1682, _d1683, _d1684,
                   _d1685, _d1686, _d1687, _d1688, _d1689, _d1690, _d1691, _d1692, _d1693, _d1694, _d1695, _d1696, _d1697, _d1698, _d1699,
                   _d1700, _d1701, _d1702, _d1703, _d1704, _d1705, _d1706, _d1707, _d1708, _d1709, _d1710}),
                    .DOBX({_d1711, _d1712, _d1713, _d1714, _d1715, _d1716, _d1717, _d1718, _d1719, _d1720, _d1721, _d1722, _d1723, _d1724,
                   _d1725, _d1726, _d1727, _d1728, _d1729, _d1730, _d1731, _d1732, _d1733, _d1734, _d1735, _d1736, _d1737, _d1738, _d1739,
                   _d1740, _d1741, _d1742, _d1743, _d1744, _d1745, _d1746, _d1747, _d1748, _d1749, _d1750}),
                    .ECC1B_ERRA({_d1751, _d1752, _d1753, _d1754}),
                    .ECC1B_ERRB({_d1755, _d1756, _d1757, _d1758}),
                    .ECC2B_ERRA({_d1759, _d1760, _d1761, _d1762}),
                    .ECC2B_ERRB({_d1763, _d1764, _d1765, _d1766}),
                    .FORW_CAS_WRAO(_d1767), .FORW_CAS_WRBO(_d1768), .FORW_CAS_BMAO(_d1769), .FORW_CAS_BMBO(_d1770), .FORW_CAS_RDAO(_d1771),
                    .FORW_CAS_RDBO(_d1772), .FORW_UADDRAO({_d1773, _d1774, _d1775, _d1776, _d1777, _d1778, _d1779, _d1780, _d1781, _d1782,
                   _d1783, _d1784, _d1785, _d1786, _d1787, _d1788}),
                    .FORW_LADDRAO({_d1789, _d1790, _d1791, _d1792, _d1793, _d1794, _d1795, _d1796, _d1797, _d1798, _d1799, _d1800, _d1801,
                   _d1802, _d1803, _d1804}),
                    .FORW_UADDRBO({_d1805, _d1806, _d1807, _d1808, _d1809, _d1810, _d1811, _d1812, _d1813, _d1814, _d1815, _d1816, _d1817,
                   _d1818, _d1819, _d1820}),
                    .FORW_LADDRBO({_d1821, _d1822, _d1823, _d1824, _d1825, _d1826, _d1827, _d1828, _d1829, _d1830, _d1831, _d1832, _d1833,
                   _d1834, _d1835, _d1836}),
                    .FORW_UA0CLKO(_d1837), .FORW_UA0ENO(_d1838), .FORW_UA0WEO(_d1839), .FORW_LA0CLKO(_d1840), .FORW_LA0ENO(_d1841),
                    .FORW_LA0WEO(_d1842), .FORW_UA1CLKO(_d1843), .FORW_UA1ENO(_d1844), .FORW_UA1WEO(_d1845), .FORW_LA1CLKO(_d1846),
                    .FORW_LA1ENO(_d1847), .FORW_LA1WEO(_d1848), .FORW_UB0CLKO(_d1849), .FORW_UB0ENO(_d1850), .FORW_UB0WEO(_d1851), .FORW_LB0CLKO(_d1852),
                    .FORW_LB0ENO(_d1853), .FORW_LB0WEO(_d1854), .FORW_UB1CLKO(_d1855), .FORW_UB1ENO(_d1856), .FORW_UB1WEO(_d1857), .FORW_LB1CLKO(_d1858),
                    .FORW_LB1ENO(_d1859), .FORW_LB1WEO(_d1860), .CLOCKA({_d1861, _d1862, _d1863, _d1864}),
                    .CLOCKB({_d1865, _d1866, _d1867, _d1868}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7115_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7116_10, na7117_9, na7119_10, na7121_9, na7123_10, na7125_9, na7126_10, na7127_9, na7128_10, na7130_9,
                   na7137_10, na7138_9, na7139_10, na7143_9, na7149_10, na7150_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7151_10, na7153_9, na7155_10, na7156_9, na7159_10,
                   na7162_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h0843c08509187a108424084040016b5ad4a4a5294a50842280421295296b421295296b0000000000),
             .INIT_01(320'h0c0210c0210c0210f020040284a54a5ad084a4000201c4d52b00000425294800000000204bc0a041),
             .INIT_02(320'hc8439c043808681c8721c8439e043c08781a063c0c021e0681c8721c8439a04340878180421e0601),
             .INIT_03(320'h0872408421c84210902108421204210842408421086010c0210a02108421090210848108681c8721),
             .INIT_04(320'ha0721c87210e4310070108421a8421a803408421cf02408421ae021084350d021084390843905021),
             .INIT_05(320'h001210e41109021086a4c0421086a109021086a4c0421086a109021086a0484392e821204210d471),
             .INIT_06(320'h884810843506021084350842d6042109421085a10c481084210c4210d421204210d451086a288435),
             .INIT_07(320'h08421a92a5cd4a5a962109021086b52c421204210d4952e6a52d4b10848108435a962109021086a1),
             .INIT_08(320'h08421a842008421a830108421a842408421a828108421c84b1254b9a94b52c421204210d6a588424),
             .INIT_09(320'h0b42188021084218d52108021086a5a9735296a58842008421ad4b108401084350c42008421a8301),
             .INIT_0A(320'h08421ae4b108401084350c421004210d401eb621004210d45d8c420a0421086a1085ac0842128421),
             .INIT_0B(320'h040390e439087211242908621404392c421004210d7258842008421a862108021086ab0872588420),
             .INIT_0C(320'h08201084290f0214841008421487010a43f095210402108521c04a908e2180721c87210e42248521),
             .INIT_0D(320'h086a108021086a0a0421086a108021086a908c21da6290a60108421484250a4090858108521f0429),
             .INIT_0E(320'h0840108435a9621004210d4710c0390e439087290c0390e439087290c0390e4390873108061a0421),
             .INIT_0F(320'ha0421086a108021086bd0a4290d4030d021084350840108435e86b00e4390e421cd4b52e6a52d4b1),
             .INIT_10(320'h80421086a108021086a148521144300e4390e421c8aa148521040390e43908722a85214843108061),
             .INIT_11(320'h0843505021084350840108435187290a43a4d52148021485210a4298842908021086a0481210a435),
             .INIT_12(320'h8842008421aaf258842008421ae4b108401084350c421004210d40d8840108435050210843508401),
             .INIT_13(320'h484208c0390e4390872950201c8721c84394a87105021084350840108435e152bc962108021086a1),
             .INIT_14(320'h6a021084a10842d086200852108431a952108021086b00a52908541080b509b46a8c66d1aa212821),
             .INIT_15(320'h5ac1805021084350842d4042109421085a10c401084210c6a54852908401084350028108421a8421),
             .INIT_16(320'h000352d4b9a96a5ad6a5294a100001a96a5cd4b52d6b5294a508000029294a5294a5094a121ca54a),
             .INIT_17(320'h0a5260c44188e214a4084e535485200a5310a5204ac21016a109725a8845c96a002021a8c2548560),
             .INIT_18(320'h0c529000018a520001200813b4d5014822148529024290002148429480010a4214a4010883100429),
             .INIT_19(320'h5803d2d4e1a97258c5208a41148229067b1a96a0cf63d4d4a1a902108421085094a4000042948000),
             .INIT_1A(320'ha833d8f425484300843c0d4b92c6294833d8d4b5067b1ea421e06a5c96314e535585200a5310a520),
             .INIT_1B(320'h0e7b1ed4254873d8d4b5067b1e84a9a94352e4b18a419ec6a5a833d8f5210f0352e4b18a419ec6a5),
             .INIT_1C(320'h2e4b1096212a439ec6a5a833d8f4254d4a1ad4b92c425884a9387810d4a1a97258c5290e7b1a96b5),
             .INIT_1D(320'h4a5294a94b5a40002008084294243de05294a5295296b480004a0210e7b1a96a1cf63d09535286b5),
             .INIT_1E(320'h3256b0852a4a5294a1244a0210a5090f7814a5294a54a5ad20001002240902489404214a121ef029),
             .INIT_1F(320'h4a400000000000948000400e94a529525292a40108528084294243de05294a5295296b4800040089),
             .INIT_20(320'h085295e4a9ca4a95f0214a5094a4000010908529022290202548061125094a400005294800002129),
             .INIT_21(320'h0a5295800040389085295e52be04294a5200010060781085294ac000200c0f0210a5295800040389),
             .INIT_22(320'h00000001000183c4812b00001eb7a94a52000100e27810a531024214ac000203d0f0214a409e2781),
             .INIT_23(320'h4a5294a1284a5284a56000100e24394ac000201c48729580004043c0d520000294a400001094a520),
             .INIT_24(320'h4b0390e4390872c0e4390e421ca52b00008003e12a5614f021ec4294a42902d29000080702a0d529),
             .INIT_25(320'h0e421c8121e0429e2501c8721c8439e04290243c08528081280f021481280e4390e421cb02909529),
             .INIT_26(320'h4800040101c8721c8439020390e43908722898200f42d0a029087b1884204852140428084280e439),
             .INIT_27(320'h4a509425294a400000000203d6878958000403814ac000201c0a5600010006d295853c0842902d29),
             .INIT_28(320'h49c240843d0a5294a4000202140721c87210e429004a18902918481087a14a481486290852900000),
             .INIT_29(320'he8529010210d4b9a97b5e8529010210d4b9af42948081086a5cd4bdaf4294802128832094612a549),
             .INIT_2A(320'hcac28084814e4214253958501085014a4280d449494294a4000203d6f6a80e4390e421cd4e120421),
             .INIT_2B(320'h4a1294802948000000004a004084352a7a14a579ed53d084a95f4212a501c8721c8439505010a129),
             .INIT_2C(320'h0e421c8442081218a45d684204a0390e439087314883120523090210c529205294a400000314a528),
             .INIT_2D(320'h0f5bd4843c4a56000101090210c5294ac0002021205390a0210252b0000940420486a7cd4e80e439),
             .INIT_2E(320'h204218a5295800040081086b14a4a14ac0002004084358a5250a5600010020421ac5292852b00008),
             .INIT_2F(320'h000094a1284a529480000000040081086b14a4a14ac00020352848108629497b10f1204ac0002021),
             .INIT_30(320'h00100404810843d0a52958000404280e4390e421c85200943120523090210f429490290c5210a520),
             .INIT_31(320'h2a4a120421e85294a94b5ac000201c490210d7a14a4f52e6a5e84a5a94b52a4e120421e85294a520),
             .INIT_32(320'h5a52a4a4b52e6a5e96a52d4a92d4b9a97a5a94b52a4b52e6a5e86a5a94b52a4b52e6a5e8625a94b5),
             .INIT_33(320'h4a4752e6a5e86a52d4a91d4b9a97a1a94b52a46100421e85294252900008010210d7a14a5694a929),
             .INIT_34(320'h20539084814e4240940120539084814e4280940108a411852938401087a14a52900008010210c7a1),
             .INIT_35(320'h0940108a411852938401087a14a5290000808401087a14a52b000080840120539084814e42409401),
             .INIT_36(320'h08401087a14a52b000080840120539084814e4240940120539084814e4240940120539084814e424),
             .INIT_37(320'h4e4240940120539084814e4240940120539084814e4240940108a411852938401087a14a52900008),
             .INIT_38(320'h084814e4240940108a411852938401087a14a5290000808401087a14a52b00008084012053908481),
             .INIT_39(320'h4a5290000808401087a14a52b000080840120539084814e4240940120539084814e4240940120539),
             .INIT_3A(320'h084814e4212052122569c8169c982949129025260a5230a5260a52baa5798e4b1c962588021087a1),
             .INIT_3B(320'h0052122569c8169c982949129025260a5230a5260a52baa5798e4b1c962588021087a14a52900008),
             .INIT_3C(320'h00450088294af31c96392c4b1004210f4294af31c96392c4b1004210f4294a52900008084814e421),
             .INIT_3D(320'h08021091212240120539084014e4240d4a1204240842448489004814e42100539084810848909120),
             .INIT_3E(320'hc962588021087a14a5798e4b1c962588021087a14a529480004a021004014e421005390903528481),
             .INIT_3F(320'h0902509425086a5090210042122424480200a72108029c8420084244848900022884414a5798e4b1),
             .INIT_40(320'h485a943520084494252b00000000094042008029c8481284a1284352848108021091212240100539),
             .INIT_41(320'h3a561481211d62048409084010f7b10c40b08c210a520001000252b0000800129024090c5280c520),
             .INIT_42(320'h0010002420484090a56000101881254ac2902423cc7bd4a5232c40908161024234a4000203110409),
             .INIT_43(320'h08429480004063c48c3c481210c789e27890c4090863c4842108529000080012102420484090a560),
             .INIT_44(320'h4f121881210c789284210a0294a40002035e24f9a843c49ca1e24090863c4f13c4862048431e2421),
             .INIT_45(320'h084214ac000203d687890f6a5c86a52842108429580004a01c4eab5386a00f1214d407024218f13c),
             .INIT_46(320'h00100e27890f6a5ad7890f6bc4863c48431e24a1084210a56000100e27890c7890c7890863c48421),
             .INIT_47(320'hef5294812102429480004000908121024204852b00008021284d529424210053102029f06294a560),
             .INIT_48(320'h4a529004291252958000400014a408ca5294a408ea5294a4010a4494a56000101080218812102423),
             .INIT_49(320'h425294800000000400014a408ca5294a408ea5294a4010a4494a5600010000529023294a529023a9),
             .INIT_4A(320'h4852b00008070210a5295800040381085294ac0000008ca4080e520184494a529480000a52900000),
             .INIT_4B(320'h0a53a4a57c4a52900008087810a53c084294a56000100e24294a52b00008071210a5294ac0002000),
             .INIT_4C(320'h0000022520000294a40000380c0529000014a520000084a52900000000014a52000101085214a520),
             .INIT_4D(320'h095210a4204813d0f03c5ac000200040528ea4080a5010a401089214853c084210a529580000a529),
             .INIT_4E(320'h094294a121284294f029580004a0002253d486250a429e86290853d0c521e042948128484a908449),
             .INIT_4F(320'h0852b00008070210a521e04294a56000100e0781c942948780086a94f0210a53c084294a52b0e521),
             .INIT_50(320'h8a4c1024034a40002000d252b0a7890c429481684a5200010001fade87810a520e04214a7810a531),
             .INIT_51(320'h000080c429e86291c4290c53b0d52138401c86a9080204ac21484001a520001018853d0c52388521),
             .INIT_52(320'h000080009d6a4384ac29e24310a5205a52900001eb4314c52900001086290c5200c5218a7114c529),
             .INIT_53(320'h1f7a1e042948fbd0f0214a47de87810a523e04294a52000100e2421e05210a5614a0294a10b5a529),
             .INIT_54(320'h020000e4390e421c80fd6a43c0a52102ca958781484690a5200000b485200000000100e24398c631),
             .INIT_55(320'h4a4000201c084290e021ca52950821e0429085290a5211a4294a12a52d6b00000424224a40000000),
             .INIT_56(320'h805204a6010a6014a52900000425094a5290000000008070210a43c0a4214ac29484290a52842d6a),
             .INIT_57(320'h085300a5084a52900009402014e529585200c0214a5205812980429805284252948000406300a461),
             .INIT_58(320'h8052bca4250c0295e521286014ac300a6010a6014a5200012804029ca52b0a401804294a40b02530),
             .INIT_59(320'h00008001300a6010c5204a6010a60148126081200052958000402014c0214c0214c0294ac0002029),
             .INIT_5A(320'h4a5610f429481684252900008001300a7294ac29804310a52902c094c0214c029024c10240842529),
             .INIT_5B(320'h024094ac00020004c02902530085300a409304090252b00008003294ac294f121485290a52a0f521),
             .INIT_5C(320'h4c0214c0294ac00020004c02902530085300a409304090252b00008001300a4094c0214c029024c1),
             .INIT_5D(320'h80530085300a5290000804021ea530087b54a6010f6a94a52b000080402980429805295800040201),
             .INIT_5E(320'hc8439e2431e24310843c0e4390e421cf0390e439087230a529000080f5bd0f12958000406300a461),
             .INIT_5F(320'h88c31e07218843100f81cf0390e4390873c4862108781c8721c8439e24310e43c4862108781c8721),
             .INIT_60(320'h8f039f06230c4618c4218f0390c4218807c0e781cf83118623086210c781c86210c403e073c0e7a1),
             .INIT_61(320'h070390e4390872932529580000240000000025018f0390e439087211078908789070390e43908722),
             .INIT_62(320'h0a5290040100822984214a509080294a4294a4012a52958000470390e43908728480294a5294a129),
             .INIT_63(320'h085294ac000201c4c52b000080712d4ac000201c4d52b00000425294800000000404200a1200a529),
             .INIT_64(320'h0010002420484090c0210a429804210a429804210a429804290a601085214c02148534084290a681),
             .INIT_65(320'h00008070310852b00008070310852b00008040214c0214c0214c0210a6010853008429804214a560),
             .INIT_66(320'h4a1294a40000000006a4eb52149ea58d4b509439ec6290a4352d6b5294a03852900008070310852b),
             .INIT_67(320'h0a52149831005284852988e230e02948c014a1214a6230e0294a120087ad0e029480214a52000008),
             .INIT_68(320'h084214a4e1404200e0210d4b92c425884a14a7010842949c2808401c042948529480004042b08121),
             .INIT_69(320'h2842108721087a8084210843d88421e84210f4410843d08421e85210853d0616b00009403010a538),
             .INIT_6A(320'h084210843d88421e84210f441087a10843d0a4210a7a0c2d60001280201c484210f4210873408421),
             .INIT_6B(320'h0f43da94200003d0f6a5080000f43da9420001280201c484210f42108734084212842108721087a8),
             .INIT_6C(320'h48429a8e2148535011394d521480294c4294812b08405a8425c96a211725a8008086a30952158000),
             .INIT_6D(320'h4d4b10a7890d4a9425284a4000240102775a903504429a8121480010a6a000429a98200c4e188e21),
             .INIT_6E(320'h2c6290262902629026290e7b1a96a1cf63d4d4a1a97258c520cf6352d419ec7a9a96a5cd4a5a9621),
             .INIT_6F(320'h8a53aad4b92c629386a00a6350a43501c152e4b18a401e86a5c96314873d8d4b50e7b1ea6a50d4b9),
             .INIT_70(320'hcf63d484280d4b92c629067b1a96a0cf63d4d4b52e6a52d4b108781a97258c529a96210f0352e4b1),
             .INIT_71(320'h8c52900435a97258c520cf6352d419ec7a908501a97258c5270f0210a0352e4b18a429067b1a96a0),
             .INIT_72(320'h00001a9725884b10952900001a97258c529000094a02102629004218a43148021eb43108781a9725),
             .INIT_73(320'h0000040301e87a1e843d4ac3808538085380f43d0f421ee1290000802829c04290a5010a52b00000),
             .INIT_74(320'h4ac00020200f0290943d480350a52b00008003890a4250f5310a529580000a529000004252948000),
             .INIT_75(320'h804210a601084294a400000000201c08521287a98a57c0a4250f529480004001c48521287a988529),
             .INIT_76(320'ha04214d0210a54a4a5294a43d4c021085244a12148521485300842148c2912449804210a60108429),
             .INIT_77(320'h48089a943548021aa5294a021ca53808529c04294e0214a58108529604250a5280842140421a0429),
             .INIT_78(320'h0a429a07a1e87a10f7a18a409085204892148bb18a52948000404340f43d0f421e9bb10d0294d029),
             .INIT_79(320'he843de862917621a0529021210b434085340f43d0f421ef431480220a681e87a1e843de862922421),
             .INIT_7A(320'h0a4b14c5340f43d0f421ef4314804148829d05210a72148029a07a1e87a10f7a18a56122681e87a1),
             .INIT_7B(320'h484a148489086290a4014f4314a4250a424484314853b0c5340f43d0f421ef431480090808908429),
             .INIT_7C(320'h8a4020a429484a148489086290a4014f4314a4250a424484314853b0c5340f43d0f421ef43148029),
             .INIT_7D(320'hef43148c218a681e87a1e843de8629204010f6210241d8c523ec6290012100121a07a1e87a10f7a1),
             .INIT_7E(320'h01e81e87a1e843daa681e87a1e843d0840108409485292862902409084290a409085340f43d0f421),
             .INIT_7F(320'h8a681e87a1e843de062900429e8629a07a1e87a10f7a18a401c56a9386b40f43d0f421ef621aa529)) 
           _a6636 ( .DOA({_d1869, _d1870, _d1871, _d1872, _d1873, _d1874, _d1875, _d1876, _d1877, _d1878, _d1879, _d1880, _d1881, _d1882,
                   _d1883, _d1884, _d1885, _d1886, _d1887, _d1888, _d1889, _d1890, _d1891, _d1892, _d1893, _d1894, _d1895, _d1896, _d1897,
                   _d1898, _d1899, _d1900, _d1901, _d1902, _d1903, na6636_36, na6636_37, na6636_38, na6636_39, na6636_40}),
                    .DOAX({_d1904, _d1905, _d1906, _d1907, _d1908, _d1909, _d1910, _d1911, _d1912, _d1913, _d1914, _d1915, _d1916, _d1917,
                   _d1918, _d1919, _d1920, _d1921, _d1922, _d1923, _d1924, _d1925, _d1926, _d1927, _d1928, _d1929, _d1930, _d1931, _d1932,
                   _d1933, _d1934, _d1935, _d1936, _d1937, _d1938, _d1939, _d1940, _d1941, _d1942, _d1943}),
                    .DOB({_d1944, _d1945, _d1946, _d1947, _d1948, _d1949, _d1950, _d1951, _d1952, _d1953, _d1954, _d1955, _d1956, _d1957,
                   _d1958, _d1959, _d1960, _d1961, _d1962, _d1963, _d1964, _d1965, _d1966, _d1967, _d1968, _d1969, _d1970, _d1971, _d1972,
                   _d1973, _d1974, _d1975, _d1976, _d1977, _d1978, _d1979, _d1980, _d1981, _d1982, _d1983}),
                    .DOBX({_d1984, _d1985, _d1986, _d1987, _d1988, _d1989, _d1990, _d1991, _d1992, _d1993, _d1994, _d1995, _d1996, _d1997,
                   _d1998, _d1999, _d2000, _d2001, _d2002, _d2003, _d2004, _d2005, _d2006, _d2007, _d2008, _d2009, _d2010, _d2011, _d2012,
                   _d2013, _d2014, _d2015, _d2016, _d2017, _d2018, _d2019, _d2020, _d2021, _d2022, _d2023}),
                    .ECC1B_ERRA({_d2024, _d2025, _d2026, _d2027}),
                    .ECC1B_ERRB({_d2028, _d2029, _d2030, _d2031}),
                    .ECC2B_ERRA({_d2032, _d2033, _d2034, _d2035}),
                    .ECC2B_ERRB({_d2036, _d2037, _d2038, _d2039}),
                    .FORW_CAS_WRAO(_d2040), .FORW_CAS_WRBO(_d2041), .FORW_CAS_BMAO(_d2042), .FORW_CAS_BMBO(_d2043), .FORW_CAS_RDAO(_d2044),
                    .FORW_CAS_RDBO(_d2045), .FORW_UADDRAO({_d2046, _d2047, _d2048, _d2049, _d2050, _d2051, _d2052, _d2053, _d2054, _d2055,
                   _d2056, _d2057, _d2058, _d2059, _d2060, _d2061}),
                    .FORW_LADDRAO({_d2062, _d2063, _d2064, _d2065, _d2066, _d2067, _d2068, _d2069, _d2070, _d2071, _d2072, _d2073, _d2074,
                   _d2075, _d2076, _d2077}),
                    .FORW_UADDRBO({_d2078, _d2079, _d2080, _d2081, _d2082, _d2083, _d2084, _d2085, _d2086, _d2087, _d2088, _d2089, _d2090,
                   _d2091, _d2092, _d2093}),
                    .FORW_LADDRBO({_d2094, _d2095, _d2096, _d2097, _d2098, _d2099, _d2100, _d2101, _d2102, _d2103, _d2104, _d2105, _d2106,
                   _d2107, _d2108, _d2109}),
                    .FORW_UA0CLKO(_d2110), .FORW_UA0ENO(_d2111), .FORW_UA0WEO(_d2112), .FORW_LA0CLKO(_d2113), .FORW_LA0ENO(_d2114),
                    .FORW_LA0WEO(_d2115), .FORW_UA1CLKO(_d2116), .FORW_UA1ENO(_d2117), .FORW_UA1WEO(_d2118), .FORW_LA1CLKO(_d2119),
                    .FORW_LA1ENO(_d2120), .FORW_LA1WEO(_d2121), .FORW_UB0CLKO(_d2122), .FORW_UB0ENO(_d2123), .FORW_UB0WEO(_d2124), .FORW_LB0CLKO(_d2125),
                    .FORW_LB0ENO(_d2126), .FORW_LB0WEO(_d2127), .FORW_UB1CLKO(_d2128), .FORW_UB1ENO(_d2129), .FORW_UB1WEO(_d2130), .FORW_LB1CLKO(_d2131),
                    .FORW_LB1ENO(_d2132), .FORW_LB1WEO(_d2133), .CLOCKA({_d2134, _d2135, _d2136, _d2137}),
                    .CLOCKB({_d2138, _d2139, _d2140, _d2141}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7168_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7169_10, na7170_9, na7172_10, na7173_9, na7174_10, na7175_9, na7177_10, na7179_9, na7180_10, na7181_9,
                   na7193_10, na7194_9, na7195_10, na7196_9, na7197_10, na7199_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7200_10, na7201_9, na7205_10, na7213_9, na7214_10,
                   na7215_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h0281f6294c5302b0280a500410084210842108421084210822108421084210842108420000000000),
             .INIT_01(320'h401e0401e0401e047c022fc421084210842108411081f10442104407884210820080005281f5294b),
             .INIT_02(320'h081e103d007a00f0bc2f081e103d007a3e003fdf001e8f800f0bc2f081e103d007a3e003c08f800f),
             .INIT_03(320'h7bfe07bdeffa108401e84210803d08421007a1084200f401e0401ee6a1e8401e00200f0200f0bc2f),
             .INIT_04(320'h03c2f0bc20785e84280f73deffbdeffa1407bdefffc007bdeff81ee7bdff401ee7bdff7bdff401ef),
             .INIT_05(320'h421ef7fd0f501ef7bfe003dcf7bfef501ef7bfe003dcf7bfef501ef7bfef7b9e17b80a03def7fde8),
             .INIT_06(320'h7a80f7bdff001ee7bdff7bdff0b9af781ee73bef7fc00001ef7fdef7fdea03def7fde87bfef43dff),
             .INIT_07(320'h7bdeffa1ef4bdef7bdef501ef7bfe97bdea03def7fd0f7a5ef7bdef7a80f7bdff4bdef501ef7bfe8),
             .INIT_08(320'h73deffbd407bdeff800f73deffbd407bdeff800f73deffa1e843de97bdef7bdea03def7fd2f7bd40),
             .INIT_09(320'h77deff80006bdeffa10f501ef7bfe87bd2f7bdef7bd407bdeffa5ef7a80f7bdff43d407bdeff800f),
             .INIT_0A(320'h7bdeffa5ef7a80f7bdff7bdea03def7fde0781ea03def7fdef7bc0003dcf7bfef7bfe1735ef03dce),
             .INIT_0B(320'h00141585810382e7bc0f03de0781e97bdea03def7fd2f7bd407bdeffbdef501ef7bfef03d2f7bd40),
             .INIT_0C(320'h0000f73d0f03de1780007b9e8781ef0bc0f781e0001ee7a1e07bc0f03de00282b0b020705cf781e0),
             .INIT_0D(320'h7bfef501ef7bfe003dcf7bfef501ef7bfef03c00721087a00f73d0e781ef720084282e789e07bc4f),
             .INIT_0E(320'h7a80f7bdff4bdea03def7fdef00141585810382f00141585810382f00141585810382f001e003dcf),
             .INIT_0F(320'h03dcf7bfef501ef7bfef6bc0f0200f001ee7bdff7a80f7bdff78100505616040e0a10f7a5ef7bdef),
             .INIT_10(320'h03d2e7a10f501ef7bfee781e07bc00505616040e0b90e781e000141585810382e439e0781ef001e0),
             .INIT_11(320'h7bdff001ee7bdff7a80f7bdff781cf03c0e4210f43daf601807bc087b9e8501ef7bfe0401e073c08),
             .INIT_12(320'h7bd407bdeffa12f7bd407bdeffa5ef7a80f7bdff7bdea03def7fd007a80f7bdff001ee7bdff7a80f),
             .INIT_13(320'h43c4f4014158581038284000a0ac2c081c1421e8001ee7bdff7a80f7bdff781084bdef501ef7bfef),
             .INIT_14(320'hf85cd7bc0f739df7bfe00010e7bdff73d0f501ef7bfe07a1087a10f109ef7e1d9c01f675ec07a1cf),
             .INIT_15(320'h1085f001ee7bdff7bdff0b9af781ee73bef7fc00035ef7fdaf439087a80f7bdff0240f73deffbdef),
             .INIT_16(320'h089ef7bdee7bdef789cf7884a1044f7bdef73def7bc4e7bc425082203c427884f109e213c4f08842),
             .INIT_17(320'h7210e021c0421ee420084390843d0f6a10f72100421e213def5c1b18016651cc05a14b42c4840842),
             .INIT_18(320'h7bc421044f78842088487f10e4210f43d0e43908021e803c0e43dc8401e0721ee4200f03c08781c8),
             .INIT_19(320'h1000f0084f7bdef7bc4f109e213c427b5af739cf631ee139ef109c2689825bc421084113de210822),
             .INIT_1A(320'h73d8c7b9a013d4043d5f7bdef7bde213dad7b9ce7b18f709eafbdef7bdef1384213c4f6884f70840),
             .INIT_1B(320'h7b5af709c013dad7b9ce7b18f7340273def7bdef789ed6bdce73d8c7b84f57def7bdef789ed6bdce),
             .INIT_1C(320'h7bdef781cf009ed6bdce73d8c7b9a0139ef13def7bde073c0212bed7bdef7bdef7bc427b5af739c2),
             .INIT_1D(320'h10842108421084110800781e2789e1fbc42108421084210822109e07b5af739cf631ee6804e7bc4f),
             .INIT_1E(320'h789ef0004f13c4f13c4f101e0789e2787ef10842108421084208840789e2789e203c0f13c4f0fde2),
             .INIT_1F(320'h1084100401101e210822101e2789e2789e27880f03c40781e2789e1fbc42108421084210822101e2),
             .INIT_20(320'h7bde2139e2709e217def7884210841101e27bde203c0203dc0101e0789e21084113de21082203c42),
             .INIT_21(320'h7bc4210822103e27bde213c42fbdef1084208840003e07bde2108411080007c0f7bc4210822103e2),
             .INIT_22(320'h080200884003d5f100421044f781ef7884208840f8bee7bc420084b10841109ef57def78802f8be0),
             .INIT_23(320'h73dc213dcf708421084208840f89e0108411081f13c021082213d5f78042089ef10841101e210842),
             .INIT_24(320'h101e1785e103c20785e17840f0884210442001ef1884f17daf7bdc2789e2008421044207c0f7544f),
             .INIT_25(320'h7840f08040fbde2f880f0bc2f081e1fbde20081f7bc400004007def10040785e17840f081c278de2),
             .INIT_26(320'h108221000f0bc2f081e1001e1785e103c2f13c0003df8501e213def109401084a03c4078040785e1),
             .INIT_27(320'h7b9ee7b8421084100401109ef02be210822103e0108411081f00842088400384213c5f781e200842),
             .INIT_28(320'h1094073c0f7884210841109e00282b0b020705e2001c0101e21280e781ef1080f13c4212c4210440),
             .INIT_29(320'h7bc42001c07bdef7bde27bc42001cf035ad13de21000e03def7bdef13de2101ee03c0e701ee009e2),
             .INIT_2A(320'h089417a82e785ea089e1128287a82f78941789ef1096210841109ef7bc40505616040e0884a039e0),
             .INIT_2B(320'h73dc21098210820080221080073c0d689ef1084e7bc4e789e2139e07880a0ac2c081c11282f5044f),
             .INIT_2C(320'h6040e0a1e05004f789ef03d4010141585810382f1380203c42501cf03c4203c4210841101e213dcf),
             .INIT_2D(320'h7bc0e03d5f108420884f501cf03c4210841109ea0b9e1505ea008421044213c0013c427884050561),
             .INIT_2E(320'h039e078842108221000e7804f1084b108411080073c02788425884208840039e013c4212c4210442),
             .INIT_2F(320'h0880f73dcf7084210820080221000e7804f1084b10841109ef7a80e781e213def57c4010841109ea),
             .INIT_30(320'h088400000e7800f788421082213c00505616040e0bc400380203c42501cf03de2101e27884258842),
             .INIT_31(320'h7884a039e07bc4210842108411081f101cf009ef1084f7b9ef6bc0273def7884a039e07bc4210842),
             .INIT_32(320'h7884f1084f7b9ef789cf7bde213dee7bde273def7884f7b9ef6bfe273def7884f7b9ef6bc0273def),
             .INIT_33(320'h1084f7b9ef789cf7bde213dee7bde273def7884a039e07bc421084210442001cf009ef109e213c42),
             .INIT_34(320'h0b9e17a82e785417880a0b9e17a82e785417880f03dc0781e21280e781ef1084210442001cf009ef),
             .INIT_35(320'h7880f03dc0781e21280e781ef10842104427a80e781ef10842104427800a0b9e17a82e785417880a),
             .INIT_36(320'h7a80e781ef10842104427800a0b9e17a82e785417880a0b9e17a82e785417880a0b9e17a82e78541),
             .INIT_37(320'h785417880a0b9e17a82e785417880a0b9e17a82e785417880f03dc0781e21280e781ef1084210442),
             .INIT_38(320'h7a82e785417880f03dc0781e21280e781ef10842104427a80e781ef10842104427800a0b9e17a82e),
             .INIT_39(320'h10842104427a80e781ef10842104427800a0b9e17a82e785417880a0b9e17a82e785417880a0b9e1),
             .INIT_3A(320'h7a82e785ea0bc4a0884f0804f0b80f13de27bc4e03c4e03c4e03c427884f139e273c4f101e0009ef),
             .INIT_3B(320'h0bc4a0884f0804f0b80f13de27bc4e03c4e03c4e03c427884f139e273c4f101e0009ef1084210442),
             .INIT_3C(320'h781ee03c0f109e273c4e789e203c0013de2109e273c4e789e203c0013de210842104427a82e785ea),
             .INIT_3D(320'h5050f5044a0880a0b9e17a82e785417bdea0bd4143d41128220282e785ea0b9e17a8287a82250440),
             .INIT_3E(320'h73c4f101e0009ef1084f139e273c4f101e0009ef1084210822109e00282e785ea0b9e1505ef7a82f),
             .INIT_3F(320'h505ef7bdef73def505ea0a1ea089411014173c2f505cf0bd4143d411282203c0f701e07884f139e2),
             .INIT_40(320'h7b80278040781e210842104010044213c00505cf0a82f7bdef7b9ef7a82f5050f5044a0880a0b9e1),
             .INIT_41(320'h7884f1004013c4010002780007bdc2788020080258842088400084210442000420080f7004f70040),
             .INIT_42(320'h088400080010002008420884f1004f109e200802789ef7bc4278802000400080210841109e212802),
             .INIT_43(320'h131621082213c5f1095f1004f00be2f8be2788027805f109c262c421044200040008001000200842),
             .INIT_44(320'h17c4f1004f00be21344c1096210841109e2f884e13d5f109eaf88027805f17c5f13c4013c02f884e),
             .INIT_45(320'h609ab10841109ef02be27bdef709cf7884e13162108221081f1384213c4857c4e10802009e017c5f),
             .INIT_46(320'h08840f8be27bdef78be27bc5f13c5f13c02f884e1304d5884208840f8be278be278be27805f109c2),
             .INIT_47(320'h7bdef100400080210822100020004000800100421044203c4f13de2789ea0bc5e03c027bfc210842),
             .INIT_48(320'h13de20380278842108221000f7880f73c4f7880f73c4f7880e009e2108420884f0000f1004000802),
             .INIT_49(320'h7884210820080221000f7880f73c4f7880f73c4f7880e009e2108420884003de203dcf13de203dcf),
             .INIT_4A(320'h100421044207c0f7bc4210822103e07bde2108411000f0880f70440781e278842108227bc4210440),
             .INIT_4B(320'h7084f1085f10842104427abef7bc5f03def1084208840f89ef108421044207c4f7bc421084110800),
             .INIT_4C(320'h1044078842089e2100411010043c421044f788420880f10842104010044f788420884f7b84e13c40),
             .INIT_4D(320'h73c4f009411004857d5f10841108007804f0880f009ee1080f03c4f13c40781c0788421082278840),
             .INIT_4E(320'h7b80f13c4e7b80f17c0210822108007884f13dee009e27bde27bc4e7bc4afbdef100427b9e2781ef),
             .INIT_4F(320'h12c421044207dcf7bc4afbdef1084208840f83ef6b80f12be173c0f17c0f7bc5f73def13c4f039e0),
             .INIT_50(320'h789ea0080210841108007084278be27bdc210042108420884003def7abef7bc40f81ef78bee7bc42),
             .INIT_51(320'h10442789e27bde213de27bc4f791e0780007bc8f03d4013c0f78000108420884f13c4f7bc427bc4f),
             .INIT_52(320'h10442001ef78940109e2f89ef70840108421044f7bdcf13c421044f7b9e27bc4073c4f789cf13c42),
             .INIT_53(320'h13deafbdef109ef57def7884f7abef7bc42fbdef1084208840f89e203c4e1084f108421084210842),
             .INIT_54(320'h10800785e17840f081ef7095f789e0009e212bef781ef008420880f100420802008840f896110842),
             .INIT_55(320'h108411081f7b84f0000c0884213c4203c0270842788427bc021084210842104407880f1084100401),
             .INIT_56(320'hfbc4010bef00bef10842104407b9ee10842104010044207dee13c00789c2109e2109ef0084210842),
             .INIT_57(320'h7805f788421084210442103ef1384213c4857dae1084010042fbc02fbc42108421082213c5f7884a),
             .INIT_58(320'hfbc42789ef57de213c4f7abef1095f78bef00bef108420884207de2708427890afb5c2108020085f),
             .INIT_59(320'h104420005f78bef7084010bef00bef1004f500401304210822103ef17de017de017de210841109e2),
             .INIT_5A(320'h1084e03dc21004210842104420005f789c2109e2fb5ef708420080217de017de2009ea0080210842),
             .INIT_5B(320'h00802108411080017de20085f7805f788027a8020084210442001c2109c217c4f13842708427384e),
             .INIT_5C(320'h17de017de2108411080017de20085f7805f788027a80200842104420005f7880217de017de2009ea),
             .INIT_5D(320'hfbc5f7805f788421044207dee7085f73def10bee7bde2108421044207de2fbc02fbc4210822103ef),
             .INIT_5E(320'h081e1f89e4f89e47805f785e17840f0fde1785e103c2200842104427bc0f57c421082213c5f7884a),
             .INIT_5F(320'h109e2fbc2f7bde200bef0fde1785e103c3f13c8f00bef0bc2f081e1f89e47841f13c8f00bef0bc2f),
             .INIT_60(320'h17de1780427884e13def17de17bdef1005f787ef0bc0213c42701ef78bef0bdef78802fbc3f785e0),
             .INIT_61(320'h07d415858103822788421082200841004011084f17d4158581038287abe27abe207de1785e103c2f),
             .INIT_62(320'h7bde20000003c0f701e0789e253dce13def788007bc421082217de1785e103c2f13dce13def13c42),
             .INIT_63(320'h03d82108411081f104421044207c41108411081f100421044078842108200802213c0003c4f7384f),
             .INIT_64(320'h08840008001000207dee009e2fb9e0789e2fb9e0789e2fbdc278bee7bc4f17dee13c5f701ec78bee),
             .INIT_65(320'h1044207de212c421044207de212c421044207def17def17def17de078bef03c5f781e2fbc0f10842),
             .INIT_66(320'h13c42108410040113c4f7804f109ef73def6bda17b1e2789ef7bc4e7bc40100421044207de212c42),
             .INIT_67(320'h7bc4f138027b44d13de21084257def109ed1344f7884257def13c4003def57def13c00108420880f),
             .INIT_68(320'h7b8027884afbd4047daf7bdee739007a00878bef7004f1095f7a808fbc0f12c421082213c025004e),
             .INIT_69(320'h03dcd6a3ee723ff0000d6a1ff7b5a8fb9c87fde07391f7b5a8fadee7201f17c4210442103ef03c5f),
             .INIT_6A(320'h0000d6a1ff7b5a8fb9c87fdee723ef6b51f5bdce403e2f8842088421001f7b9ad47dce43fe0735ef),
             .INIT_6B(320'h7bdef10942089ef7bc42508227bdef10942088421001f7b9ad47dce43fe0735ef03dcd6a3ee723ff),
             .INIT_6C(320'h43dc8421ee439080210e4210f43da843dc8401087884f7bd706c600599473016852d0b1210210822),
             .INIT_6D(320'h139ef78be27bde210842108411090fe21c8421e87a1c84010f401e072100781c843c0f021c0421ee),
             .INIT_6E(320'h7bde2789e2789e2789e27b5af739cf631ee139ef7bdef7bc4f6b5ee739ec63dc273def73def7bdef),
             .INIT_6F(320'h7884e13def7bde213c4f689c2709e2009ef7bdef78800781cf7bdef13dad7b9ce7b18f709cf7bdef),
             .INIT_70(320'h631ee13d5f7bdef7bde27b5af739cf631ee139ef7a1ef7bdef4abef7bdef7bc4243de857def7bdef),
             .INIT_71(320'h7bc42001c27bdef7bc4f6b5ee739ec63dc27abef7bdef7bc4257d0f57def7bdef789e27b5af739cf),
             .INIT_72(320'h0044f7bdef7bc0e780421044f7bdef7bc4210442109e0789e2001cf789ef1000f781ef42bef7bdef),
             .INIT_73(320'h08022103ea0ac2c081c11095f7bc5f7bc5f785e17840f080421044203c02fbdc278bef0084210401),
             .INIT_74(320'h10841109e057def73dc11000f0084210442003e27bdcf7044f00842108227bc42104407884210820),
             .INIT_75(320'h03c007880f001e210841004011081f6bdee7b8227885f7bdcf70442108221001f13dee7b82278042),
             .INIT_76(320'hfbc0f17de0789ef7bdce739c1101e003c4f13c4f13c4f13c407800f13c02789e203c007880f001e2),
             .INIT_77(320'h101e273def13c0f709ef17dcf3bc5f781e2fbc0f17de078bef03de2fb9e07bc5f78002fbc02fbde2),
             .INIT_78(320'h789e2fbc2f0bc20785e0788027bc4013c4f13def788421082213c1f785e17840f0bdef57def17def),
             .INIT_79(320'h081e1781e27bdeafbde203c4e7a95f7bc5f785e17840f0bc0f1000f00bef0bc2f081e1781e2009cf),
             .INIT_7A(320'h789cf13c5f785e17840f0bc0f101c0138027804e009e013802fbc2f0bc20785e07884a00bef0bc2f),
             .INIT_7B(320'h7b9e81280273de27880f13def13dcf40940139ef13c4f03c5f785e17840f0bc0f100020000273de2),
             .INIT_7C(320'h7880f009e27b9e81280273de27880f13def13dcf40940139ef13c4f03c5f785e17840f0bc0f101e2),
             .INIT_7D(320'h0bc0f1380f78bef0bc2f081e1781e2780007bdea009ef7bc4f7bde20004000040fbc2f0bc20785e0),
             .INIT_7E(320'h00bea0ac2c081c178bef0bc2f081e1780007a9e27bde2701e20080273de2788027bc5f785e17840f),
             .INIT_7F(320'h78bef0bc2f081e1781e2001e27bde2fbc2f0bc20785e078800709e213c5f505616040e0bdee13de2)) 
           _a6637 ( .DOA({_d2142, _d2143, _d2144, _d2145, _d2146, _d2147, _d2148, _d2149, _d2150, _d2151, _d2152, _d2153, _d2154, _d2155,
                   _d2156, _d2157, _d2158, _d2159, _d2160, _d2161, _d2162, _d2163, _d2164, _d2165, _d2166, _d2167, _d2168, _d2169, _d2170,
                   _d2171, _d2172, _d2173, _d2174, _d2175, _d2176, na6637_36, na6637_37, na6637_38, na6637_39, na6637_40}),
                    .DOAX({_d2177, _d2178, _d2179, _d2180, _d2181, _d2182, _d2183, _d2184, _d2185, _d2186, _d2187, _d2188, _d2189, _d2190,
                   _d2191, _d2192, _d2193, _d2194, _d2195, _d2196, _d2197, _d2198, _d2199, _d2200, _d2201, _d2202, _d2203, _d2204, _d2205,
                   _d2206, _d2207, _d2208, _d2209, _d2210, _d2211, _d2212, _d2213, _d2214, _d2215, _d2216}),
                    .DOB({_d2217, _d2218, _d2219, _d2220, _d2221, _d2222, _d2223, _d2224, _d2225, _d2226, _d2227, _d2228, _d2229, _d2230,
                   _d2231, _d2232, _d2233, _d2234, _d2235, _d2236, _d2237, _d2238, _d2239, _d2240, _d2241, _d2242, _d2243, _d2244, _d2245,
                   _d2246, _d2247, _d2248, _d2249, _d2250, _d2251, _d2252, _d2253, _d2254, _d2255, _d2256}),
                    .DOBX({_d2257, _d2258, _d2259, _d2260, _d2261, _d2262, _d2263, _d2264, _d2265, _d2266, _d2267, _d2268, _d2269, _d2270,
                   _d2271, _d2272, _d2273, _d2274, _d2275, _d2276, _d2277, _d2278, _d2279, _d2280, _d2281, _d2282, _d2283, _d2284, _d2285,
                   _d2286, _d2287, _d2288, _d2289, _d2290, _d2291, _d2292, _d2293, _d2294, _d2295, _d2296}),
                    .ECC1B_ERRA({_d2297, _d2298, _d2299, _d2300}),
                    .ECC1B_ERRB({_d2301, _d2302, _d2303, _d2304}),
                    .ECC2B_ERRA({_d2305, _d2306, _d2307, _d2308}),
                    .ECC2B_ERRB({_d2309, _d2310, _d2311, _d2312}),
                    .FORW_CAS_WRAO(_d2313), .FORW_CAS_WRBO(_d2314), .FORW_CAS_BMAO(_d2315), .FORW_CAS_BMBO(_d2316), .FORW_CAS_RDAO(_d2317),
                    .FORW_CAS_RDBO(_d2318), .FORW_UADDRAO({_d2319, _d2320, _d2321, _d2322, _d2323, _d2324, _d2325, _d2326, _d2327, _d2328,
                   _d2329, _d2330, _d2331, _d2332, _d2333, _d2334}),
                    .FORW_LADDRAO({_d2335, _d2336, _d2337, _d2338, _d2339, _d2340, _d2341, _d2342, _d2343, _d2344, _d2345, _d2346, _d2347,
                   _d2348, _d2349, _d2350}),
                    .FORW_UADDRBO({_d2351, _d2352, _d2353, _d2354, _d2355, _d2356, _d2357, _d2358, _d2359, _d2360, _d2361, _d2362, _d2363,
                   _d2364, _d2365, _d2366}),
                    .FORW_LADDRBO({_d2367, _d2368, _d2369, _d2370, _d2371, _d2372, _d2373, _d2374, _d2375, _d2376, _d2377, _d2378, _d2379,
                   _d2380, _d2381, _d2382}),
                    .FORW_UA0CLKO(_d2383), .FORW_UA0ENO(_d2384), .FORW_UA0WEO(_d2385), .FORW_LA0CLKO(_d2386), .FORW_LA0ENO(_d2387),
                    .FORW_LA0WEO(_d2388), .FORW_UA1CLKO(_d2389), .FORW_UA1ENO(_d2390), .FORW_UA1WEO(_d2391), .FORW_LA1CLKO(_d2392),
                    .FORW_LA1ENO(_d2393), .FORW_LA1WEO(_d2394), .FORW_UB0CLKO(_d2395), .FORW_UB0ENO(_d2396), .FORW_UB0WEO(_d2397), .FORW_LB0CLKO(_d2398),
                    .FORW_LB0ENO(_d2399), .FORW_LB0WEO(_d2400), .FORW_UB1CLKO(_d2401), .FORW_UB1ENO(_d2402), .FORW_UB1WEO(_d2403), .FORW_LB1CLKO(_d2404),
                    .FORW_LB1ENO(_d2405), .FORW_LB1WEO(_d2406), .CLOCKA({_d2407, _d2408, _d2409, _d2410}),
                    .CLOCKB({_d2411, _d2412, _d2413, _d2414}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7223_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7225_10, na7226_9, na7227_10, na7229_9, na7230_10, na7231_9, na7236_10, na7237_9, na7238_10, na7239_9,
                   na7241_10, na7242_9, na7243_10, na7244_9, na7246_10, na7247_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7248_10, na7249_9, na7251_10, na7252_9, na7253_10,
                   na7254_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h0100d211a05b00c07005402001000443214c700443214c7320ffbbc8c1ee6b16a398a10000000010),
             .INIT_01(320'ha5400a341fa4400a542587e19c5ed5a4e49406000700960141002007310b5400000004200152017c),
             .INIT_02(320'h05e80a0304061140001804b808028c05126a001d28408893140001801e00c011005323e800888820),
             .INIT_03(320'h823e902210fe39486400c729048198e52190531ca40a084402820000711483401042200c11400018),
             .INIT_04(320'h0500006001400067818002200fa214fbc1902208f943902214fb0004401f404004411f4421f07408),
             .INIT_05(320'h03d8887de004008853f080008803e006008853f080008803e006008853e003f0013d8080110a7c05),
             .INIT_06(320'h002804429fac0004401f4421f2000058090443e887e016891027d1087c00a0110a7dc2443ee1a21f),
             .INIT_07(320'h02214fbe107c2088400404008853f080060e0110a7df083e1044200100804429f8400104008853ef),
             .INIT_08(320'h02200f801102214f838002200f801002214f92a002208fd0097c20f84110800c0e0110a7e1001408),
             .INIT_09(320'h87d10ff42e02204fa88006408853ef841f0822100081902214fc200080a04429f7800902214fa500),
             .INIT_0A(320'h02214fbd00102a04429f00020e8110a7dc0fbc0068110a7c1f0e001e8008803e8843f00000b01208),
             .INIT_0B(320'h2168000300200000101c000007000f800c0e8110a7de80140902214f800404408853ee001f000c09),
             .INIT_0C(320'h021200229c03bc02038500114e01de0100ef0080254004538077804000000d00006008a000020380),
             .INIT_0D(320'h803e002408853e108008803e002408853e0038207b1af0b3200228fe01d00300078020f808077804),
             .INIT_0E(320'h082a04429f84000e8110a7c180528000300a300801280003009f00405280003009201806000a8008),
             .INIT_0F(320'h28008803e006408853ee7a00403980024004401f003a04429f701cca0000c033c039f083e1044200),
             .INIT_10(320'h08000451c204408853ef403800001ca0000c0170001cf4038041280003003900073d00e000002000),
             .INIT_11(320'h4429f210004401f001804429f001e40200f439e1439ece01600a00403c4804008853e8071c07a00e),
             .INIT_12(320'h0101802214fbdf000c0802214fbd00102804429f00020e0110a7def000804429f264004401f00180),
             .INIT_13(320'hc00000d28000300e301cc51140001806380e6001a20004401f003804429f7030f7a00504008853e0),
             .INIT_14(320'hfe40002c048221f443e40ae004409f8430002008853f807218451e003c8478ea3e800398fa003be0),
             .INIT_15(320'h5a80d000004401f4421fa000058090443e887c015811027e10c3f84001804429f0008002200fa210),
             .INIT_16(320'h040108420f8421043a10439e080200842107c210821d0821cf040000399c7438ea71d8e3b94039ac),
             .INIT_17(320'h7a08ff6dfddbc0f2708003d8a7858e7b3807b19003c007908f00de3e800368fa002be05000b50100),
             .INIT_18(320'h0158a802001b150003800010f229e123b6f63d0403c2803bcf605e8221dd7b02f4118ef3bbb775ec),
             .INIT_19(320'h0704e069fb841c80818e4b1ca6396c738018410d6801f6420513c0f03c0f001ca40600800cc54010),
             .INIT_1A(320'h435a02fde06001d0000d0420e4040c639c00c2086b400fb000e82107202063f9a7878e7f1807f090),
             .INIT_1B(320'h73809fe9e0639c0442086b407fbc0c8439083901031ce00610435a007d800541083901031ce01a10),
             .INIT_1C(320'h8390a6812e031ce02210435a03fde06420ec420e421a03b80c781a004202841c80818c7380a8411a),
             .INIT_1D(320'ha419c7358b50600830090061c77200c83148338e6b16a0c010430007380a8410d6813f7819083b10),
             .INIT_1E(320'h071cd00380e0380e0380e4401a71dca0000c520ce39ac5a830041800701c0701ce8034e3b8c03018),
             .INIT_1F(320'h5aa00000008000c540106001c0701c0701c07200083990069c77300403148338e6b16a0c0106001c),
             .INIT_20(320'h0300c7bc447f0285440c0318b50600801cc0200c0380ca3800621c10200c5aa008000c5401003988),
             .INIT_21(320'h0018a08010600380300c7878a681806283000380200210400c5040007000074008018a0801060238),
             .INIT_22(320'h0000000380000016014100200fbc202315000380ab0200018b031e0504000701f044040310c2b23f),
             .INIT_23(320'h234046388d0218c5a82000380ab10050400070016000a0801060015000300400062a00801cc42d50),
             .INIT_24(320'h6100040380b200c00100e02a002d410020c001d9071e1e7400f81fc8310ce01418001c0740e0198e),
             .INIT_25(320'he013404190c810c0b3200201c01380e810c6303502191e2181504086319d00100e032405008d020c),
             .INIT_26(320'h0c000e03200201c06a006140040380b2000580080b8000100ce03e15bc18601e0a03880038d00100),
             .INIT_27(320'h721a46810c5aa00000000701f783aa08000e00a15040007009028200418003d1c7878507d0c2016a),
             .INIT_28(320'h63c190009f6318b50600830008c01804014c018cc05e1fe40c780a0007ec631a06396c7814180200),
             .INIT_29(320'hfb18c0640404201843defb18c2640024201f7d8c661a0202100421ef7d8c661c40384f401c8021c8),
             .INIT_2A(320'h03c0d000a020000270007838000220830050281063c0a406008301f0879d2030060158071e0e8004),
             .INIT_2B(320'h2340863c0b54000000104301100110863ec631effa30ff81187bc01263240601405580c03a002388),
             .INIT_2C(320'h202e800017001806301f7a40865400600808b00c63c3fa018f004000b18c2018a40600801c76390d),
             .INIT_2D(320'h07def000156282000380040000b18c5040007000a800004000c3141002086003c6038f0700d00180),
             .INIT_2E(320'h6000f6318a08000e038000d4c631e050400070000004a6318f0282000380280015318c781410001c),
             .INIT_2F(320'h0400e4348d0218b5400000000e038001d4c631e05040007010802800018c603e1025805040007000),
             .INIT_30(320'h00380a20000001f6318a080106001ce0080e0264031980bc3f2018f040000fd8c6600c72d8f02830),
             .INIT_31(320'h851e0e001dfb39c7358b5040083019620000fbec631f083e107fc1e84190821e0e0001fb18c5a830),
             .INIT_32(320'h7538ec71f083e107ba10242107c20f843ee840d0861f083e107ffee84190831f083e107fc0e841d0),
             .INIT_33(320'h631f8c3f187ff18263047e30fc63ffc60d8c21e088005fb18c62d418001c02000ebbece71cce3a1c),
             .INIT_34(320'ha8100001806000907900a810000180200080788e081e270a0c782a003fec631418020c030002ffec),
             .INIT_35(320'h0788e081e270a8c780a0043ec631418001c000a003fec631410020c00100a8280001808000907900),
             .INIT_36(320'h002a0043ec631410020c001002028000380800190790020100003806001907900201000038020019),
             .INIT_37(320'h0000907900a010000180e000907900a010000180c00090788e081e270b0c782a004fec631418001c),
             .INIT_38(320'h00380c00190788e081e270b8c780a0053ec631418001c000a004fec631410020c00100a028000180),
             .INIT_39(320'h631418001c002a0053ec631410020c00100202800038000019079002010000380e00190790020100),
             .INIT_3A(320'h0038060000a03806e1e8041e403c386020c0618f0c18f0e18f0c18f161eebbd167c2b8a3417253ec),
             .INIT_3B(320'ha83806e1e8041e403c3c6028c0718f0d18f0f18f0d18f161eebbd167c2b8a3418253ec631418020c),
             .INIT_3C(320'h7040f1385863dd67a2af85313c006787d8c63dd37a24f847104804487d8c629018020c0038060000),
             .INIT_3D(320'h0640003380e600020100003a0e0018042002801000004e0298c038040000a8300001800003c04310),
             .INIT_3E(320'h7c2989f0033c3ec631ee9bd127c23883002243ec631480c01043000401a0a0000280000001080180),
             .INIT_3F(320'h0000370dc10021002000a800047018c000102000064180001100004e0298c3820789c2e31eeb3d15),
             .INIT_40(320'h7100c701887040862d4100000002086000802414000800b86e08010801800640003380e608028100),
             .INIT_41(320'h061ffc0180787f86078c0010107dff02c8f43c0f0283000380231410001c021840300e2018e00188),
             .INIT_42(320'h00380e30006038c0a82004180fd180c3ff8e300f77fe10218f0fe8c0d1e8a300050600830177808c),
             .INIT_43(320'h7800a0c010603f163c05601800afac2b3ac02a8c0017163c0f001418001c06180a30286058c02820),
             .INIT_44(320'h665805418002dac781e07b80a406008301eab1eff001563d004b08c0056162581601586000bab1e0),
             .INIT_45(320'h03c00504000701f781ac07f187ab180ade07800a080104300163d1e787cf0358f27980e30015e581),
             .INIT_46(320'h00380ab1ac07e10421ac07d01601596000bab1e0781e00282000380ab1ac027ac02aac0017163c0f),
             .INIT_47(320'h0fc0860181a300a0c000e028c0018123000605410001c0018e6040c73000401002382c700085a820),
             .INIT_48(320'h6008c23c280216a08000e01a00300e211802308ed91802308f0a0085a820041800a000fe181e300f),
             .INIT_49(320'h7310b5400000000e03a00300e111802308ee91802308f0a0085a820003802800c038246008c23bc4),
             .INIT_4A(320'h601410001c044004118a08000e00a10208c504008000e0328e00188704087218b540100018a80200),
             .INIT_4B(320'h7f10e4714162d418001c0032081189081846282000380ea00462d410001c045002118b504000700c),
             .INIT_4C(320'h80200031500400c78200800080018a80200031500400e6216a800000020043150041800bd0fe0180),
             .INIT_4D(320'h7890c03c19601ef0741d404000700070d8e0300e131c00300e1010060194000004316a08010031e0),
             .INIT_4E(320'h03c246398f130046540a08000c7000031ee603ef0a1c4f85047349f02080280802608f03c4860000),
             .INIT_4F(320'h781410001c01400a0180282806282000380887a07bc24600310500465420c018d002806118e03f00),
             .INIT_50(320'h4b0008300050600830007938f0f12c001fc4300c5a83000380003e1083a06018088408031200018b),
             .INIT_51(320'h8020c07dccf852c7a1cc0258ef87800010177c3c0000c63801e001c0283004180fb99f0a58f43980),
             .INIT_52(320'h8020c0001f7700143c3c8b0007f10c02d4180200f85e86258a8020003d2c021807a580431e96218a),
             .INIT_53(320'h78fe0a818063c5f0640c031e1f83a060180a818062830041808b00080100071e823e1183dcd62d41),
             .INIT_54(320'h8300c40280603300301f7e01c0738003c6c78380e001c028300400e6015000000041800b200e77df),
             .INIT_55(320'h506008700d0018003410073148018ca000c0318fa21f00001183dcd62d41802007300062a0000000),
             .INIT_56(320'h6818c620201b0a062d4180200711a04316a800000020c01400e000c0301ce3c887c0000460f7358b),
             .INIT_57(320'h00d89031ac5a901802086002063c1c7878f0040fe1190051884806c6818d62d480c010603e5031e0),
             .INIT_58(320'hc818f770100440c7bb80402a063c0903220fb2a0628300410c0740c7838f0f1e0e81fc2320083105),
             .INIT_59(320'h8001c041940322001d9c622201328067180001807816a08000e002067419634066400c504008301c),
             .INIT_5A(320'he01ef07dfc4500d62d418020c04194031e0e3c3c400007f08c8010c470026000c430006300d62d41),
             .INIT_5B(320'h6300b50400070086300c03114001980300c0008c02d410020c001e0e3df4e1580a3f847f10f03f0f),
             .INIT_5C(320'h630066400c50400070186700c8310400d880320c0028c02d410001c041940310c470126000c43000),
             .INIT_5D(320'h6019401598031418001c03000fa184003e84300007e0862d410001c0300c4008c6018a08000e0200),
             .INIT_5E(320'h059800b0216b02102a1c402002027001100800809400f0a9018001c07de10558a08010603e4031e0),
             .INIT_5F(320'hf3c3e410008081e802140110080080df018604205610804004065008b02120158604205110804004),
             .INIT_60(320'hff1807278f0f00fe6040e708006040e30040020c0393d787a07fc82076040008207580c4004601c9),
             .INIT_61(320'h01000002005b0080216a0801002a000000082180f910080080930000018c0032c85100800808c000),
             .INIT_62(320'h4000ce008043820789c2231cc0000060080030800018a08000e1100002009a00060000600006390c),
             .INIT_63(320'h0000c5040007019601410001c00580504000700960141002007310b5400000000e00080818000180),
             .INIT_64(320'h003808300c6010c040004b18c6000b6338c6000a6318ce800c632a00318c670006619d0040063320),
             .INIT_65(320'h0001c0140b781410001c0140b781410001c0700c6301c6700c62410633a0fb19400b0c8011862820),
             .INIT_66(320'h6390c5aa0000000003c0fbddf43e107c20078600fbc0d0b010823d0823cc7fd6a0001c0740b78141),
             .INIT_67(320'h0118463fde73d8c6048cf3faf03400601cf63181233ef0340060188003e101400638a05a83004000),
             .INIT_68(320'h0005c031e0e800d020001420f421c03bc020318000bc063c1900320003c0601480c0106002f03100),
             .INIT_69(320'h05202743e27c3f50a0227c29f589f0f89f087dc113e1f709f0f81427c01f2fd010020860300f0190),
             .INIT_6A(320'h0a0227c29f589f0f89f087c027c3ee13e1f0284f803e5fa0200031c280096004f87c4f843e00000b),
             .INIT_6B(320'h07cdf73c100401f3fdcf0401007cff73c100031c280196004f87c4f843f00000b05202743e27c3e5),
             .INIT_6C(320'he05e833c0fe3d060000f629e1639ece01ec6400f001e423c0378fa000da3e800af814002d4040010),
             .INIT_6D(320'h44200120a80420462d494060007000021ea33c2676dec361e1401dd7b0dc779ec33bceee9fddbc0f),
             .INIT_6E(320'h4082c730a873088730687380b8410d6815f6421b841c81058e70050821ad007ec842107c20884001),
             .INIT_6F(320'h5310ff420e42d4c787ce7b01e7a0dea00108390b53002702107216a639c04c2086b408fb210e420e),
             .INIT_70(320'h6803f600180420e4082c738078410d680df6421083e1044200781a0841c85a9888400f004108390b),
             .INIT_71(320'h5a988405fc841c83998e70050821ad007ec00100841c81058f0500001010839020b02c738028410d),
             .INIT_72(320'h00200841c8334057018a80200841c80818a80204430007306cc11e10300367060fbc40783a0841c8),
             .INIT_73(320'h000106030c0400003680e3c00021940218c6020000150015418001c0380c8000c432200314100000),
             .INIT_74(320'h504000700005400789806300e6b1410001c020a8001e2a018e6b16a080100018a802007310b54000),
             .INIT_75(320'hc0000c32000030c5060000000830090000f1100c0f15d001e22018a0c000e01194000f1100c7358b),
             .INIT_76(320'h803f06301f831cd62d88202006300029980601806018060194000996384c0300c40008030000230c),
             .INIT_77(320'h651cc840246382e2320c614000a19d0048c0802461401230008608cc0080c119500418c8038c020c),
             .INIT_78(320'h5b10c8a00403019001cb5b22c0618560180603e1a31480c0106002d40080e0174003e10141066410),
             .INIT_79(320'h0280072d6c07c208820ca398f064000418d40080600680396b6502e0b3280100c0760072d6c03000),
             .INIT_7A(320'h631f962d9d40080602c00396b661f5c3e787330f661d0c3e180a0040300f001cb5b1e0431280100c),
             .INIT_7B(320'h6bc446038c0018ccb18e67c2c635e2230106000c6658ef319d40080600440396b6210c1630c0016c),
             .INIT_7C(320'h5b38e0b00c6bc446038c001accb18e67c2d635e2230106000d6658ef359d40080602040396b6200c),
             .INIT_7D(320'h0396b63c20731080100c0280072d6c0010107c206301f0b980f86ac01184a51838a0040301e201cb),
             .INIT_7E(320'ha01080100c06080233080100c05f00001010000c0200c78d6c8332c0016c9320c0019c400806021c),
             .INIT_7F(320'h331080100c01e8072d6c805ccf856c0200403000c01cb5b1027f88c787dc400806035407c0ff418c)) 
           _a6638 ( .DOA({_d2415, _d2416, _d2417, _d2418, _d2419, _d2420, _d2421, _d2422, _d2423, _d2424, _d2425, _d2426, _d2427, _d2428,
                   _d2429, _d2430, _d2431, _d2432, _d2433, _d2434, _d2435, _d2436, _d2437, _d2438, _d2439, _d2440, _d2441, _d2442, _d2443,
                   _d2444, _d2445, _d2446, _d2447, _d2448, _d2449, na6638_36, na6638_37, na6638_38, na6638_39, na6638_40}),
                    .DOAX({_d2450, _d2451, _d2452, _d2453, _d2454, _d2455, _d2456, _d2457, _d2458, _d2459, _d2460, _d2461, _d2462, _d2463,
                   _d2464, _d2465, _d2466, _d2467, _d2468, _d2469, _d2470, _d2471, _d2472, _d2473, _d2474, _d2475, _d2476, _d2477, _d2478,
                   _d2479, _d2480, _d2481, _d2482, _d2483, _d2484, _d2485, _d2486, _d2487, _d2488, _d2489}),
                    .DOB({_d2490, _d2491, _d2492, _d2493, _d2494, _d2495, _d2496, _d2497, _d2498, _d2499, _d2500, _d2501, _d2502, _d2503,
                   _d2504, _d2505, _d2506, _d2507, _d2508, _d2509, _d2510, _d2511, _d2512, _d2513, _d2514, _d2515, _d2516, _d2517, _d2518,
                   _d2519, _d2520, _d2521, _d2522, _d2523, _d2524, _d2525, _d2526, _d2527, _d2528, _d2529}),
                    .DOBX({_d2530, _d2531, _d2532, _d2533, _d2534, _d2535, _d2536, _d2537, _d2538, _d2539, _d2540, _d2541, _d2542, _d2543,
                   _d2544, _d2545, _d2546, _d2547, _d2548, _d2549, _d2550, _d2551, _d2552, _d2553, _d2554, _d2555, _d2556, _d2557, _d2558,
                   _d2559, _d2560, _d2561, _d2562, _d2563, _d2564, _d2565, _d2566, _d2567, _d2568, _d2569}),
                    .ECC1B_ERRA({_d2570, _d2571, _d2572, _d2573}),
                    .ECC1B_ERRB({_d2574, _d2575, _d2576, _d2577}),
                    .ECC2B_ERRA({_d2578, _d2579, _d2580, _d2581}),
                    .ECC2B_ERRB({_d2582, _d2583, _d2584, _d2585}),
                    .FORW_CAS_WRAO(_d2586), .FORW_CAS_WRBO(_d2587), .FORW_CAS_BMAO(_d2588), .FORW_CAS_BMBO(_d2589), .FORW_CAS_RDAO(_d2590),
                    .FORW_CAS_RDBO(_d2591), .FORW_UADDRAO({_d2592, _d2593, _d2594, _d2595, _d2596, _d2597, _d2598, _d2599, _d2600, _d2601,
                   _d2602, _d2603, _d2604, _d2605, _d2606, _d2607}),
                    .FORW_LADDRAO({_d2608, _d2609, _d2610, _d2611, _d2612, _d2613, _d2614, _d2615, _d2616, _d2617, _d2618, _d2619, _d2620,
                   _d2621, _d2622, _d2623}),
                    .FORW_UADDRBO({_d2624, _d2625, _d2626, _d2627, _d2628, _d2629, _d2630, _d2631, _d2632, _d2633, _d2634, _d2635, _d2636,
                   _d2637, _d2638, _d2639}),
                    .FORW_LADDRBO({_d2640, _d2641, _d2642, _d2643, _d2644, _d2645, _d2646, _d2647, _d2648, _d2649, _d2650, _d2651, _d2652,
                   _d2653, _d2654, _d2655}),
                    .FORW_UA0CLKO(_d2656), .FORW_UA0ENO(_d2657), .FORW_UA0WEO(_d2658), .FORW_LA0CLKO(_d2659), .FORW_LA0ENO(_d2660),
                    .FORW_LA0WEO(_d2661), .FORW_UA1CLKO(_d2662), .FORW_UA1ENO(_d2663), .FORW_UA1WEO(_d2664), .FORW_LA1CLKO(_d2665),
                    .FORW_LA1ENO(_d2666), .FORW_LA1WEO(_d2667), .FORW_UB0CLKO(_d2668), .FORW_UB0ENO(_d2669), .FORW_UB0WEO(_d2670), .FORW_LB0CLKO(_d2671),
                    .FORW_LB0ENO(_d2672), .FORW_LB0WEO(_d2673), .FORW_UB1CLKO(_d2674), .FORW_UB1ENO(_d2675), .FORW_UB1WEO(_d2676), .FORW_LB1CLKO(_d2677),
                    .FORW_LB1ENO(_d2678), .FORW_LB1WEO(_d2679), .CLOCKA({_d2680, _d2681, _d2682, _d2683}),
                    .CLOCKB({_d2684, _d2685, _d2686, _d2687}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7264_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7267_10, na7268_9, na7269_10, na7270_9, na7272_10, na7273_9, na7274_10, na7275_9, na7280_10, na7283_9,
                   na7284_10, na7285_9, na7287_10, na7288_9, na7289_10, na7302_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7303_10, na7304_9, na7306_10, na7307_9, na7308_10,
                   na7309_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h4651f000000741a46518d8348c0800000000002108421086bef7bdef7bdeffffffffff0000000005),
             .INIT_01(320'he2800e241fe0800e70008fffef7bdef7bffffc000801e06000f80000000007c0000003c101f00003),
             .INIT_02(320'h004a0801c803a6401003004802826304ec07481600814b82c40100300460b029007320b8014d0080),
             .INIT_03(320'hf17f9003c5fb9b32d00773665882ee6ccae061cd997402b40028c000341372c000390003a2401003),
             .INIT_04(320'h1100400c033003ef0240003d5f83d4ff80e003c5f9c1a003d4fd00007abfa3000078bf078bff3000),
             .INIT_05(320'hf78a0f7fc006400f53e1d8000f57e006400f53e3e8000f57e006c00f53e00022006800f001ea7f7e),
             .INIT_06(320'h0020007a9fc280007abf07a7fa00000029307be0f7ea00001ea7c1ea7c00a001ea7e9e07bf4f03df),
             .INIT_07(320'h003d4ff400000000000002800f53e0000005801ea7fa00000000000001c007a9f0000003c00f53fd),
             .INIT_08(320'h003d5f801f003d4f8180003d5f8001003d4f8920003c5fe03de800000000000003001ea7c0000008),
             .INIT_09(320'hf7c1efe400003d4ff68006000f53fd00000000000001c003d4f8000003c007a9fe801f003d4f9c20),
             .INIT_0A(320'h003d4f80000022007a9f000009001ea7c4838000a001ea7f670051d70000f57e0f4ff80000005260),
             .INIT_0B(320'h128802006031c00009014084812000000005801ea7c000000d003d4f800003800f53e14000000010),
             .INIT_0C(320'h4136000261407e0120b9000130a03f00901f804845c0004c280fc02424484100400c064000012028),
             .INIT_0D(320'hf57e005c00f53e1d8000f57e006400f53e240408efbbe07ae0002600a0000785ee8340f80481fc02),
             .INIT_0E(320'h0020007a9f000008801ea7f2145080200603ac0245880200603a80245c80200603a8014782810000),
             .INIT_0F(320'h98000f57e001c00f53e200902476414580007abf0014007a9f123af20080180eb077a00000000000),
             .INIT_10(320'h7000004fa000400f53e01202818904200801810d003a01202811c802006043000e80480a04243c28),
             .INIT_11(320'h07a9f0680007abf0030007a9f0a0024091cf77c0f00000a048009140001e07800f53e3f0c480091d),
             .INIT_12(320'h00010003d4ff40000012003d4f80000026007a9f00000a001ea7fc0002c007a9ff040007abf002c0),
             .INIT_13(320'he800af2880200604c01de858401003025c0ef43e9dc0007abf0016007a9f103bd0000003c00f53e0),
             .INIT_14(320'hf840000014983df07be3003a007a9f003a000800f53f5077bd04fa000000000000000000000077e0),
             .INIT_15(320'h003f40480007abf07a7fd80000029307be0f7fa00001ea7c00e83b40038007a9f30300003d5f83d3),
             .INIT_16(320'h0000000000000000000000000f80000000000000000000000007c010000000000000000001300000),
             .INIT_17(320'h07fe41f803f7800ff8ffffbfef83e007fc007fc1ff8000000000000000000000007fe0f001ef083e),
             .INIT_18(320'h00000f80000001f0083e003f8ffbe0f83c0f03ff0fc1f00040f001ff840207800ffc411807e00c1e),
             .INIT_19(320'h068000001f0000000000000000000000000000000000700000000000000000000087c00000007c00),
             .INIT_1A(320'h0000001c000001a0001f000000000000000000000000038000f80000000007800000000000000001),
             .INIT_1B(320'h000003800000000000000000038000003e00000000000000000000001c0006c00000000000000000),
             .INIT_1C(320'h000000000000000000000000001c0000000000000000000000002a00000000000000000000000000),
             .INIT_1D(320'h0000000000007c00840300180000e01000000000000000f801084000000000000000070000000000),
             .INIT_1E(320'h7802100001004010040106c00000008036000000000000003e004200802008020f80000000d07c00),
             .INIT_1F(320'h003e0000000000007c01080401004008020080a00041500000002e0a800000000000000f80108200),
             .INIT_20(320'h0000000000000000680000000007c0000000000000300000180040000000003e00000007c0000000),
             .INIT_21(320'h0000007c01082200000000000980000003e00400b828000000003e008019054000000007c01082e0),
             .INIT_22(320'h000000040007c1e00000f8000380000001f00400c01800000018000003e00800703c00000a0e01e7),
             .INIT_23(320'h0000000000000000001f00400d0018003e00801c0030007c000001e0601f00000003e0000000001f),
             .INIT_24(320'h00ac0a828005803b02a0a001400001f0021003b40000003800380000000008001f002006c00f4000),
             .INIT_25(320'ha003802000d80009837605414006e0d80005801e0001773c18078000441fb02a0a001705400a0000),
             .INIT_26(320'h0f8020825605414007200d2c0a82800e4010f4000010002c01004e00840a004205000000019b02a0),
             .INIT_27(320'h0000000000003e000000080070038007c01003e0003e0080000001f00420078000001901c0008000),
             .INIT_28(320'h000170000700000007c00840026c1a06800c8000080000500000120000e0002800000000001f0000),
             .INIT_29(320'h3800000c0000000002e038000114000000801c0000ce0000004001701c000144e000e6e009c00000),
             .INIT_2A(320'h0001c00280f8000383e000300002a0000160012000000087c00840700017e8340e003b0000070000),
             .INIT_2B(320'h000000000007c00000010841500000000e00000038000f800000300001fd0681e007a0002c00141f),
             .INIT_2C(320'h0000100008040000004705c11010200000007c0000400a00000240000000a0000087c00000000000),
             .INIT_2D(320'h01c000001d0001f004000440000000003e008000880600640068000f802108006000000800108000),
             .INIT_2E(320'h380000000007c01003800000000000003e00801f00000000000001f00400080000000000000f8020),
             .INIT_2F(320'h00000000000000007c0000001002a00000000000003e008000000800000007ce005400003e008000),
             .INIT_30(320'h00400dfd00000070000007c010800420080180030000100000a80000240001c0005000000000003e),
             .INIT_31(320'h00020780003800000000007c00841801800000e0000000000007c000000000000a8000380000003e),
             .INIT_32(320'h000000002000000f040000000080000032100000000200000007fe100000000200000007c0100000),
             .INIT_33(320'h0000000000f00000000000000000000000000000f00013800000001f004106400004e00000000000),
             .INIT_34(320'h300a0002c02801e00080400a00030028000000c2000c02000000380000e000001f002103800080e0),
             .INIT_35(320'h000c2000c02000000220000e000001f002000260000e000000f802100000200a0002802801c00040),
             .INIT_36(320'h000e0000e000000f802100000c80a0001002801000040d80a0001402801200080e80a00018028014),
             .INIT_37(320'h3000500040780a0003e02800700080880a00002028009000c2000c020000000a0000e000001f0020),
             .INIT_38(320'h002a02801d000c2000c02000000340000e000001f002000380000e000000f802100000680a0003a0),
             .INIT_39(320'h00001f002000200000e000000f802100000100a0002203001900040200a0002602801b00080300a0),
             .INIT_3A(320'h002c03000030000700060000600000004000800000001000000000000000000000000005000000e0),
             .INIT_3B(320'he8000280060000600000004000800000001000000000000000000000000002c00000e000001f0021),
             .INIT_3C(320'h1800b01c00000000000000000f800001c000000000000000001000001c0000021f0021001a030000),
             .INIT_3D(320'h0780006c00a8080000a0001e02801700000180020001f003203806028000980a0000a0000400700a),
             .INIT_3E(320'h0000003400000e000000000000000004000000e0000010f801084000038028000600c005000003e0),
             .INIT_3F(320'h01400000000000004400800006800702012014000040500013000100014050c00580e00000000000),
             .INIT_40(320'h00300060020800000000f8000000210800002805000200000000000001a0030000240018080700a0),
             .INIT_41(320'he001f05c0000017002600000001c0000060003800003e0040068000f802003800080000600006001),
             .INIT_42(320'h004007000b002600001f004200181d003e088000000e0000000026000800c0000007c008400001c0),
             .INIT_43(320'h000000f80108019000130380000300d81c0001e00001a0000000001f0020040004000d001200001f),
             .INIT_44(320'h00c0001000001e00000000000087c008400980000000d0000070120000140580a0000a00000a8000),
             .INIT_45(320'h00000003e008007003a001c0000000000000000007c010840d078000000001c00000201000003410),
             .INIT_46(320'h004000028001c00002a001c16000160000008000000000001f004002832000320003400000500000),
             .INIT_47(320'h01c0001c00580000f80100100024002800e00000f80200000000000000004c80008000048000001f),
             .INIT_48(320'h00000104000000007c01003a0000000000000020f800000041000000001f00420000000240028000),
             .INIT_49(320'h0000007c000000100280000000000000020f800000041000000001f00400c80000000000000083e0),
             .INIT_4A(320'h00000f8020060000000007c010034000000003e000000c000006001000000000007c0000000f8000),
             .INIT_4B(320'h000000001d00001f00200024000012000000001f004009800000000f80200540000000003e008002),
             .INIT_4C(320'hf8000f001f0000007be000300c0000f80000001f0000000000f8000000000001f004200000000001),
             .INIT_4D(320'h000024000c0180005c19003e00800000000c002000000c00410000802000000080000007c000001e),
             .INIT_4E(320'h0000000000009000380007c0100000d0000003e0001003810000007020009000002c000000012060),
             .INIT_4F(320'h00000f80200100000000300000001f0040040140000000017a034000200000009000000000040008),
             .INIT_50(320'h403e058000007c008400f00000034000000004000003e00400078e00002000000080000004000000),
             .INIT_51(320'hf802100100381000000002001d8048e800006c024040700900120000003e00420020070200000000),
             .INIT_52(320'ha8021003c70001500000480000000100001f00003800802000f80004010002001020004002802000),
             .INIT_53(320'h000e020000000070140000000380c000000380000003e02920c8001f80000801f0014a5294948009),
             .INIT_54(320'h084025012048008007c7000180000800000002e0020404003e000000201f0000000420b80c000000),
             .INIT_55(320'h026a094405000214090a00000000293810002631f80121851294800000116800008100003e000000),
             .INIT_56(320'hb8013003600024000001f00000000000000f800000149004000050700000423e0028414294a52529),
             .INIT_57(320'h000090000000021f0021081a0078000000004c000000103c00b800070000000010f8010801200000),
             .INIT_58(320'h10000000000200000000001200000a001a0200800003e0042101c00f000000000680000002050012),
             .INIT_59(320'hf00200641b000600001c00080003600641f014000000007c010000001c040200307c00003e008400),
             .INIT_5A(320'h0000041c0000c0000001f002104c15003c000000f0000000000830007c0005c00a83e00000000001),
             .INIT_5B(320'h88000003e00800a03000680140040b00140f82a000000f8021003800000005800000000000000000),
             .INIT_5C(320'h0280000400003e008002010002800d0000400040f81a000000f802001808001200400202000303e0),
             .INIT_5D(320'hf80020001900001f00200100038005000e0000c001c0000000f80200000040000f800007c0100040),
             .INIT_5E(320'h019c020380103800003368180600cd055a06018032c0100042e802001c000700007c010801a00000),
             .INIT_5F(320'h0840184400f804108630031a06018033c1c07000001cd0300c019e0d83805801f070000062d0300c),
             .INIT_60(320'h09e20e8021004200f8020a620078020882b90171074010802101fe0105b1003e0104417440f883c0),
             .INIT_61(320'h1eb20c02e0058000800007c00003e000000108400f9a0601803d0000032000080101a0601803c801),
             .INIT_62(320'h00000080401000010020000000000000000000a00000007c0105f40c02e006400000000000000000),
             .INIT_63(320'h05000003e00801b06000f802007418003e00801e06000f80000000007c0000001000000000000000),
             .INIT_64(320'h0040040007000c00600010080c800200060d000200060d00001036000001070000000400280000a0),
             .INIT_65(320'hf80200300000000f80200400000000f802005004054030540305400102a00041c01c00b80400001f),
             .INIT_66(320'h00000003e0000000801c3801f0000000000003403800000000000000000307c00f802002c0000000),
             .INIT_67(320'h04000074600001000200000000240000000040008000002c0004006000e005800004080003e00010),
             .INIT_68(320'h00000000005800f07400000000000000000003e0000000000f00220e8060000010f8010800003400),
             .INIT_69(320'h07fc0007e0007fa00000007fff8001f8001fffe00003ff8001f83e00041f07c21f0021082c01801b),
             .INIT_6A(320'h00000007fff8001f8001fffe0007ff0003f07c00083e0f843e008210000ff80000fc000fbf900000),
             .INIT_6B(320'h01c070001f0000701c0007c0001c070001f0082100005f80000fc000fbef0000007fc0007e0007f1),
             .INIT_6C(320'hf001fff800f03ff37ffeffbe0f801ff001ff07fe000000000000000000000001ff83c007bc20f800),
             .INIT_6D(320'h00000002200000000001087c0107c007f3effc1f0781ef83e0f800307be000c1ef844117843f7800),
             .INIT_6E(320'h000000000000000000000000000000000070001f00000000000000000000000e0000000000000000),
             .INIT_6F(320'h0001d0000000000000000000000000080600000000300000000000000000000000000038000f8000),
             .INIT_70(320'h000070000b0000000000000000000000007000000000000000003800000000000000000740000000),
             .INIT_71(320'h000002000000000000000000000000000e00012000000000000180002c0000000000000000000000),
             .INIT_72(320'h00000000000000000000f80000000000000f80210840000000000000000000400383800016000000),
             .INIT_73(320'h000010814c02c0b00180000060000b0000d601605800a00c01f002000200d00000010000000f8000),
             .INIT_74(320'h003e00800006800001e00040000000f80200038000000680010000007c0000000f80000000007c00),
             .INIT_75(320'hd00042036001000007c0000000841300000044000001500000880000f80100016000000440008000),
             .INIT_76(320'h103ec0041f6016b5ac00002c0054000300c0300c0300c030170000b02c0000000c80015034000500),
             .INIT_77(320'h001800000c000006000001c110000f0000090000050000030028000581c00000b0000040000d8180),
             .INIT_78(320'h601601581506002b8020602c00201a0000c018e0000010f80108007b02a0a0053078e00480002400),
             .INIT_79(320'h00f4008180d9c0020000e300017c0f0301db02a0c00790040c07000003f60541800b000818018000),
             .INIT_7A(320'h5802b03012b02a0c007c0040c0524202c20a9805302c7008e0bd81506003d8020600007033605418),
             .INIT_7B(320'h00000000e0001805818c01c0c000000000a0000c02c020300eb02a0c009d0040c047800464000180),
             .INIT_7C(320'h6004000180000010000000180580ac01c0c00000080030000c02c0203007b02a0c009e0040c02980),
             .INIT_7D(320'h0040c03800603760541801400081800800001c0030027030013800002c0002c000581506004f8020),
             .INIT_7E(320'h10256054180146060276054180142030000000000000008580b0300001805814002818b02a0c00a0),
             .INIT_7F(320'h6015605418018802018048180381806d815060061802060180e81800000fb02a0c00a301c0000000)) 
           _a6639 ( .DOA({_d2688, _d2689, _d2690, _d2691, _d2692, _d2693, _d2694, _d2695, _d2696, _d2697, _d2698, _d2699, _d2700, _d2701,
                   _d2702, _d2703, _d2704, _d2705, _d2706, _d2707, _d2708, _d2709, _d2710, _d2711, _d2712, _d2713, _d2714, _d2715, _d2716,
                   _d2717, _d2718, _d2719, _d2720, _d2721, _d2722, na6639_36, na6639_37, na6639_38, na6639_39, na6639_40}),
                    .DOAX({_d2723, _d2724, _d2725, _d2726, _d2727, _d2728, _d2729, _d2730, _d2731, _d2732, _d2733, _d2734, _d2735, _d2736,
                   _d2737, _d2738, _d2739, _d2740, _d2741, _d2742, _d2743, _d2744, _d2745, _d2746, _d2747, _d2748, _d2749, _d2750, _d2751,
                   _d2752, _d2753, _d2754, _d2755, _d2756, _d2757, _d2758, _d2759, _d2760, _d2761, _d2762}),
                    .DOB({_d2763, _d2764, _d2765, _d2766, _d2767, _d2768, _d2769, _d2770, _d2771, _d2772, _d2773, _d2774, _d2775, _d2776,
                   _d2777, _d2778, _d2779, _d2780, _d2781, _d2782, _d2783, _d2784, _d2785, _d2786, _d2787, _d2788, _d2789, _d2790, _d2791,
                   _d2792, _d2793, _d2794, _d2795, _d2796, _d2797, _d2798, _d2799, _d2800, _d2801, _d2802}),
                    .DOBX({_d2803, _d2804, _d2805, _d2806, _d2807, _d2808, _d2809, _d2810, _d2811, _d2812, _d2813, _d2814, _d2815, _d2816,
                   _d2817, _d2818, _d2819, _d2820, _d2821, _d2822, _d2823, _d2824, _d2825, _d2826, _d2827, _d2828, _d2829, _d2830, _d2831,
                   _d2832, _d2833, _d2834, _d2835, _d2836, _d2837, _d2838, _d2839, _d2840, _d2841, _d2842}),
                    .ECC1B_ERRA({_d2843, _d2844, _d2845, _d2846}),
                    .ECC1B_ERRB({_d2847, _d2848, _d2849, _d2850}),
                    .ECC2B_ERRA({_d2851, _d2852, _d2853, _d2854}),
                    .ECC2B_ERRB({_d2855, _d2856, _d2857, _d2858}),
                    .FORW_CAS_WRAO(_d2859), .FORW_CAS_WRBO(_d2860), .FORW_CAS_BMAO(_d2861), .FORW_CAS_BMBO(_d2862), .FORW_CAS_RDAO(_d2863),
                    .FORW_CAS_RDBO(_d2864), .FORW_UADDRAO({_d2865, _d2866, _d2867, _d2868, _d2869, _d2870, _d2871, _d2872, _d2873, _d2874,
                   _d2875, _d2876, _d2877, _d2878, _d2879, _d2880}),
                    .FORW_LADDRAO({_d2881, _d2882, _d2883, _d2884, _d2885, _d2886, _d2887, _d2888, _d2889, _d2890, _d2891, _d2892, _d2893,
                   _d2894, _d2895, _d2896}),
                    .FORW_UADDRBO({_d2897, _d2898, _d2899, _d2900, _d2901, _d2902, _d2903, _d2904, _d2905, _d2906, _d2907, _d2908, _d2909,
                   _d2910, _d2911, _d2912}),
                    .FORW_LADDRBO({_d2913, _d2914, _d2915, _d2916, _d2917, _d2918, _d2919, _d2920, _d2921, _d2922, _d2923, _d2924, _d2925,
                   _d2926, _d2927, _d2928}),
                    .FORW_UA0CLKO(_d2929), .FORW_UA0ENO(_d2930), .FORW_UA0WEO(_d2931), .FORW_LA0CLKO(_d2932), .FORW_LA0ENO(_d2933),
                    .FORW_LA0WEO(_d2934), .FORW_UA1CLKO(_d2935), .FORW_UA1ENO(_d2936), .FORW_UA1WEO(_d2937), .FORW_LA1CLKO(_d2938),
                    .FORW_LA1ENO(_d2939), .FORW_LA1WEO(_d2940), .FORW_UB0CLKO(_d2941), .FORW_UB0ENO(_d2942), .FORW_UB0WEO(_d2943), .FORW_LB0CLKO(_d2944),
                    .FORW_LB0ENO(_d2945), .FORW_LB0WEO(_d2946), .FORW_UB1CLKO(_d2947), .FORW_UB1ENO(_d2948), .FORW_UB1WEO(_d2949), .FORW_LB1CLKO(_d2950),
                    .FORW_LB1ENO(_d2951), .FORW_LB1WEO(_d2952), .CLOCKA({_d2953, _d2954, _d2955, _d2956}),
                    .CLOCKB({_d2957, _d2958, _d2959, _d2960}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7330_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7331_10, na7332_9, na7333_10, na7336_9, na7337_10, na7338_9, na7340_10, na7341_9, na7342_10, na7349_9,
                   na7350_10, na7351_9, na7352_10, na7355_9, na7356_10, na7357_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7358_10, na7364_9, na7365_10, na7366_9, na7368_10,
                   na7369_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'he3d8f6338c6718fe3d8c7b1ec6318ce318c6338ce318c6318ffbdef7fdff7fdff7bfef6318c6318c),
             .INIT_01(320'h7b18c7b38f7b18c7bd8c73dad6b5ad6b7ad6b7cc6318f63d8c7b18ce318ce3d8c6719c6798f6318c),
             .INIT_02(320'h6338c631ec63d8c6318c6318c671ec63dfc6718f6358ffb18c6318c6338c631ec63dec6318f7b18c),
             .INIT_03(320'h7b9ece31ee7bdef7b38e7fdef671cf7bdec639ff7bd9c7b18c7b18c67d8f7b58ce3dac63d9c6318c),
             .INIT_04(320'h6318c6718c6318f7b38c631ed7b1fc7bd8d631eefbd8c631ec7f18c63daf7b78c63dcf63ddf7b58c),
             .INIT_05(320'h7bdcc7bdec6718c7b1ec6318c7b5ec6318c7b1ec6318c7b7ec6318c7b1ec6318c67d8c6318fe3def),
             .INIT_06(320'h6318c63d8f6b18ce3daf63d8f6b18c6318c63fec7bd8c6318f63d8fe3d8c6318f63d8f63dec7b1ef),
             .INIT_07(320'h631ec7bdbc6358c6b18c6318c7b1ed6318c6318f63ded631ac6358ce318c63d8f6b18c6318c7b3ef),
             .INIT_08(320'h631ed7b18d631ec7f18c671ed7b18c631fc7b19c631ee7b98f7b59c6f19d6718ce318f63dbc6319c),
             .INIT_09(320'h7bd8f7b58ce31ec7bdec6358c7b1ef6b19d631ac6318d633ec7b58c631bc63d8f7b19d631ec7b58c),
             .INIT_0A(320'h631ec7b18c631ac63d8f6318c6b18f67d8c6318c6b18f63d8c6318c6b18c7b5ec7b1ece318c6318c),
             .INIT_0B(320'h6318c6318c6318c6318c6318c6319c6718c6b18f63d8c6718d631ec7b38c6358c7b1ec6319c6318d),
             .INIT_0C(320'h631ac631ece31ec6318d6318f6318f6318c7b18c6358c67d8c63d8c6318ce318c6718c6318c6319c),
             .INIT_0D(320'h7b5ec6318c7b1ec6318c7b5ec6318c7b1ec6318c7bdef67dac631ec631ac63d8f7b18c7b18c63d8c),
             .INIT_0E(320'h6318c63d8f6b18ce318f63d9c6358c6318c6318c6358c6318c6318c6358c6318c6318c6358c6b18c),
             .INIT_0F(320'h6318c7b5fc6318c7b1ec6b18c67dac6318c63faf6319c63d8f631ed6318c6318c63ded631ace358c),
             .INIT_10(320'h6318ce3dec6338c7b1ec6318c6318d6318c6318c631ec6318c6358c6338c6318c7b38c6338c6758c),
             .INIT_11(320'he3d8f6f58c63faf631ac67d8f6318c6318f7bdec7b19c6319c6318fe318f6358c7b1ec7b18c6318f),
             .INIT_12(320'h6319d671fc7bd8ce319d631ec7b18c631ac63d8fe319c6b18f63fec631ac63d8f6318c63dafe31ac),
             .INIT_13(320'h7f18c7b18c6338c6318ffb18c6718c6338c7bd9f6359c63dafe31ac63d8fe31efe338c6378c7b1ec),
             .INIT_14(320'hfb18c6718c671efe3dfd633ec67d8fe31fc6378c7b1fc63defe3dec6758c6319c6338c6338c63dec),
             .INIT_15(320'h631efe318ce3fafe3d8f6f18c6338c67decfbd9c6338f63d8c7b3ef6319c63f8f6719c631ed7b1ec),
             .INIT_16(320'he318c6758c6b18ce31ac6719c7f19c671ace358c6319d6718ce3d9c6338c6718c6719c6318c6318c),
             .INIT_17(320'he3dfc67d8cfbd8c7fd8f7bdeffb1fc63dec67decfbd8c6b38c6718c6318c6718c63dec7b18f7b18f),
             .INIT_18(320'h6338c7b18c6338f6318f631ef7bdec7b1ec7f1efe3d9f6318c7b18f7b18c63d9c7bf8c6718f6318f),
             .INIT_19(320'he318c6318fe318c6719c6719c6338c6318ce318c6338c6318c6718c6318c6319c631ec6318c63d8c),
             .INIT_1A(320'he318c6319c6318c6338e6319c6338c6718c6338c6318ce319c7718ce319c63f8c6718c6338c6718c),
             .INIT_1B(320'h6338c6319c6319c6319c6338c6719c671fc6338c6318c6318c6318c6719c63b8c6318c6718c6318c),
             .INIT_1C(320'h6318ce318ce319c6318ce318ce318c6718c6718c6338c6338c631dc6319c6318ce318ce338c6318c),
             .INIT_1D(320'h6318c6718c633ec6318de318c671ec7319c6318ce318ce3d9c6318ce318ce319c6318ce318ce319c),
             .INIT_1E(320'h6318c6318c6318c6318c6318c6318c631ec6318c6318c6718f6318c6318c6318c6318c6319f63d9c),
             .INIT_1F(320'h631ece318ce318c63d9c6319c6718c6718c6318c6338ce338c6338c7b18ce318c6318c63d9c6318c),
             .INIT_20(320'h6318ce318c6338c67d8c6718c631ece318c6318c671ec631df6318ce318c671ec6338c63f8c6319c),
             .INIT_21(320'h6338c67d8ce31fc6338c6718cfb19c6338f6718ce31fc6338c671ece319c63f8c6718c63f8c631fc),
             .INIT_22(320'he338ce319c63d8f6338cfb18ce319c6338f6718cfb1fc6318ce319c633ece318c63d8c6718c7b3ec),
             .INIT_23(320'h6338c6718ce319c6319f6718c7b1cf631ec6318f679ec63d8c6718f77d9fe338ce33ec6718c6338f),
             .INIT_24(320'he318c6318c6718c6318c6318c6318c7b18c631ed6318c63d9c6319c6719c6719c7b38c63d8c7f19c),
             .INIT_25(320'h6318ce318c7338cfb3ace319c6318c7318c6318e6318deb18d6398c6318d6318c6318c6318c6b18c),
             .INIT_26(320'he3d8c633ac6318c6338c6378c6718c6338c63d9c631ac6378c6318c6319c6719c6f19d6338d6318c),
             .INIT_27(320'h6318c6318c631ec6318c6318c671cc63d8c631dc631ec6318fe318f6338c63f8c6318ee318c6338c),
             .INIT_28(320'h6319c6318c6318c631ec6318c6f18c6318c6318c6318ce318c671ace338ce338c6718c6318c7b18c),
             .INIT_29(320'h6318c6358c6318c633ec6338c6758ce319c6338c671ace318c6338f6318c6718e631ac6318c6318c),
             .INIT_2A(320'he319c633ac6718ce319c6318c6318c6318c6319c6318c631ec6318c6318c6318c6718c6718c6719c),
             .INIT_2B(320'he319c6319ce3d9c6338c6339c6338c6718c6719c6718c7b18c633ec6718c6318c6718c6318c6318c),
             .INIT_2C(320'h6b18d6718c6318ce318c63d8c633ac6b1ac6318c6318c6f18c6318c6718c6f18c631ec6338c6718c),
             .INIT_2D(320'h6718c6718fe318f6718c6758c6338c633ec6319c6b1bc6358ce318cfb18c6718c6719c6318c6b1bc),
             .INIT_2E(320'h6b38c6319c63d8c671ac6338c6318ce31ec6718d6718ce318c6718f6718ce318c6718c6718cfb18c),
             .INIT_2F(320'h6318c6318c6318c63d8c6318c631ac6318c6318c633ec6318d631ac6318c63d8c63d8ce31ece318c),
             .INIT_30(320'h6319c631ac6318ce318ce3f8c6338d6b1ac6b19d6719c6319c6318c6758c6318c6318ce318c6318f),
             .INIT_31(320'h6318c6718ce318ce318c631fc6318f6358ce318c6338d631bc63d8ceb18d6718c6718c6338c6319f),
             .INIT_32(320'he319c6338d671acfb1ac6758c6378c6f1eceb38d6318d631bc63deceb18de318d671ac63f8c6b19d),
             .INIT_33(320'h6318de31ac7b1bc6358ce378ceb38c6f38d6319c6b18c6318c6318cfb18ce338ce338c6738c6718c),
             .INIT_34(320'h631ac631ac6b18d6318c631ac633ac6b38c6738c6318c6718c671bc6719c6338c7b38c6318c6319c),
             .INIT_35(320'h6318c6318c6318c631ac6318c6318c7b18c631ac6318c6338c7b18c6318c631ac631ac6b18d6318c),
             .INIT_36(320'h631ac6338c6318c7b38c6318c6b1ac631ac6f19d6719c6b3ac631bc6f19d6719c6b3ac631ac6b18d),
             .INIT_37(320'heb18de318c6f1ac6718c6b38d6338ceb1ac631aceb18d6338c6318c6718c631ac6319c6318c7b18c),
             .INIT_38(320'h6338c6f18c6338c6338c6718c6338c6338c6718c7b38c6338c6718c6338c7b38c6319c6b1bc6318c),
             .INIT_39(320'h6319c7b18c6318c6318c6318c7b18c6718c6f1ac6319c6b18ce318c6b3ac6319c6b18c6718c6b3ac),
             .INIT_3A(320'h6318ceb18ce318c6338d6318d6318c6718c6318c6318c6318c6318c6b18c6318c6318c6318c6318c),
             .INIT_3B(320'h6b38c6319d6318d6338c6338ce338ce319c6318c6318c6b18c6718c6318ce318c6318ce318c7b18c),
             .INIT_3C(320'h6318c6318ce318ce338c6718c6b38c6318c6319c6318ce318c6318c6338c6318c7b18ce318c6b38c),
             .INIT_3D(320'h6358c6358c6b38c671ac631aceb38d6358c6718c6318de31ac6319c6b18c6b1ace318ce318c6358c),
             .INIT_3E(320'h6318c6358c6318c6718c6318c6338c6358c6338c6718c63d9c6338c631ac6b18c6b1ac6359d633ac),
             .INIT_3F(320'h6358c6318c631ac6358ceb18c6b18d6318d6358c6358d6318d6319d631ac6718c6318c6318c6318c),
             .INIT_40(320'h631ec63d8c6338ce338c7f18c6338c6318c6358d631ac6318c6318de71ace358c6358c6b18c6b1ac),
             .INIT_41(320'h7b19f6359c6318d631ac6718c6318c6318c631ec6318f6338c6319c7b19c6358c6318c77d8c73d9c),
             .INIT_42(320'h6318c6f18d633ace318f6319c6378f671ec6b18ce318ce318c633ac6319c6b18ce31fc6718c633ac),
             .INIT_43(320'h6318c67d8ce318f6318f6718c671fc7b1ec6318c6318f6318c6318c7b18c6359c6b18d631ac6318f),
             .INIT_44(320'h63d8c6318c631ece319c6318c631fc6319c7b38c6319f6338c7b18c6718f67d8f6318c6318c7b18c),
             .INIT_45(320'he318ce31ec6318c631cc671ac631ac6318c6718c63f8c6718f63d8c6318c67d8ce318c6318c63d8f),
             .INIT_46(320'h6338c7f1cc6319c633cc6318e6318f6318cfb18ce318ce338f6318cfb3cc633cc631ec6318f6338c),
             .INIT_47(320'h6718c6338c6719c63f8c6318c6319c6318c6319c7b38c6718c6318c6318c6718c6318c6319c6318f),
             .INIT_48(320'h6318c6318c6318c63d8c6318c6318c6718ce318c7b18c6319c6318c6718fe318c6319c6318ce318c),
             .INIT_49(320'h6718c63d8c6338c6318c6319c6318c6318cfb18c6318c6738c6318fe318c6318c6319c6718c631ec),
             .INIT_4A(320'h6319c7f18c63d8c6318c63d8c631ec6319c633ec6318c7b18c73d8c6318c6319ce3d8c6718c7b18c),
             .INIT_4B(320'h6b18c6318f6319c7b19c631ece318fe319c6738f6338cfb18c6318c7b38ce3d8c6719c671ec6318c),
             .INIT_4C(320'hff18c7319f6318c639ece318c6318cfb18ce338f6338ce319c7b18c6318c6319f6718ce318d6318c),
             .INIT_4D(320'h6319c6319c6318ce3d8fe31ec6718c6338c7b18c6318e7b18ce318c6338ce718c6318c63d9c6318f),
             .INIT_4E(320'h6318c6319c6318c67d8ce3d8ce338c7b38ce31fc6318c6318c6319c6718cfb18c6318c6318c6318c),
             .INIT_4F(320'h6318cff18c63d8c6718c7b38c6318f6338c7b1fc6318c631fc63d8ce3d8c6318f6319c6718c6338c),
             .INIT_50(320'h631ec6319c631ece318c7b18c631ec6318c6318c6718fe318c63d8c633ece318c7f19c671ec6319c),
             .INIT_51(320'h7b18c6718c6338c6318c6318c7b18c7b18ce3d8c6318c6318c6318ce318f6718c6338c6318c6319c),
             .INIT_52(320'h7b19c631ec6318c6718c7b18ce319c6719c7b18c631ace318c7f18c6358c6338c6b19c6318c6318c),
             .INIT_53(320'h6318c7318c6318c6398c6318c631cc6318c7318c6318f6318c7b38c6718ce318f6319c6318c6318c),
             .INIT_54(320'h6318c6b1bc6b18d633ece318f6318c6338c671ec6318c6318f6718ce338f6318c6319c7b1ac6318c),
             .INIT_55(320'h631ece338f6338c6718d6718c6718c6318c6338c7b18c6718c6319c6718c7f18ce318ce31ece318c),
             .INIT_56(320'hf318d673cc671cc6318c7b38c6318c6318c7b18c6738c67d8ce318c6318c631fce319c6318c6318c),
             .INIT_57(320'h6338ee318c6318c7b18c631cc63d8c6318c6398c6338c6358c7318c7318c6318c63d8c6318e6318c),
             .INIT_58(320'h7318c6319ce7b8ce319ce31cc6318e631cc631cce339fe339c6398c7b39c6318c7718c6718c6b38e),
             .INIT_59(320'h7f18c6319f631dc6318c631cce31ec6339f6358ce738c63f8c631cc6798c6798ce3f8c631ec6319c),
             .INIT_5A(320'h6318d6718ce318ce318cfb18ce319f673ec6338c7b18ce318c6718ce3d9c63f8ce33eceb39c6738c),
             .INIT_5B(320'he318ce33fc6318ce7f8c6318f6718fe318c7b19c6718c7b18c631fc6319c63d8c6318c6719c6718d),
             .INIT_5C(320'h24d0023e9c203ece718ce3d9c6319f6718f6338cfb18c6338cfb19c6318f6319c63f9c63f8ce31ec),
             .INIT_5D(320'h310872108621084ff08421c842108721084e70e4210842108439084e7c84390843108421c8424160),
             .INIT_5E(320'h210a4390e4310e4e7087290a42908521ca4ef0a4214842108439084e708421c8421c8421086e7084),
             .INIT_5F(320'h84210b948439084a006100c20ad2b4a5697a4e1084271a6719c6338f70e42908721c84210e5e7485),
             .INIT_60(320'ha1cbc9820ca619845d0427da024c08a0083cf3ed05f80a1084210e4a10e5210e4a000018403ac270),
             .INIT_61(320'h249b068324846102419024c9c06060020108138080a34ec334e0510a7060a426c85fb00c1b4e0794),
             .INIT_62(320'h600846418c06088220040721ce3008000844020c0000004e10848308c22084418000080030484210),
             .INIT_63(320'h0190cc0060e7193a6e987909860c97442746001762c1c1931ce300400c886601804314e0218a7010),
             .INIT_64(320'h0000420390a111006f000000018000e0304ff1802000453300a60d8a328800a942401f613dc600e0),
             .INIT_65(320'hd910422d80620845911442c880418cbf38c06e1460e0c04c148580c07044e7186814003009804297),
             .INIT_66(320'ha520ca127cc229060017441070103844400872202031083190200110110401d045800842d04c400c),
             .INIT_67(320'h6139440f1040310a708ca708c8680886008e5184e5184c4900c410001104258984501c05097a738c),
             .INIT_68(320'h613944031058310a7c8ca708c8600886008e51e4e5184c4103c41003b29c2329c02e180221861794),
             .INIT_69(320'h84e7080060000630000000063193001830038c7ce738f7f00c7f06c2329f23e9c1a2180227861397),
             .INIT_6A(320'ha228461373db31c190185de6ce71e32101324c80461647d38700000000031800000c0084e7084210),
             .INIT_6B(320'he728060203272806020027e8060208c439703010451971b01003c1484c7002288c4d6ca207042167),
             .INIT_6C(320'h1801318f9c7d0fba1e679dff059307fa203981ef442b48311ca730002200040139a2e882e6422d10),
             .INIT_6D(320'h2179c210e421084210842107000068a4c73b8e9304c071c0e05d39c62c7405217dd308a1e0819e08),
             .INIT_6E(320'h2139c2108421084210842939d21085210a4210872139c2108421084210842139c210a42148429084),
             .INIT_6F(320'hce39f21084214a4210842139c2108421084210852939c21484210a5214842939c290852108439084),
             .INIT_70(320'h212842108721280000000829184211842a421085212a000400002d4a5294ad6908c21084a98c6319),
             .INIT_71(320'h0d41484188822140c488052984121025084402e0a4298a611440f8801d94a439c600880428421084),
             .INIT_72(320'h800000229c0500820200dc280a521483010ba000c228085180202040121ce3004403e80424000214),
             .INIT_73(320'h842100424240802853c8c010300183c400a10244101024400818098861105529020174210881c010),
             .INIT_74(320'h000600000000c00000400000000000180040006000000940108401084e10842109c0008401084e10),
             .INIT_75(320'h080000002000000000600000000003000000080000003000001000000c0000003000000080000000),
             .INIT_76(320'h1806000c030000000000000400040000000000000000000001000000000000000080000002000000),
             .INIT_77(320'h0000000000000000000000c0100003000001800000c0000040080001004000002000001000010000),
             .INIT_78(320'h00000188020080010000000000000100000000000000000c0000003100401000200c000080000800),
             .INIT_79(320'h000400000000000100000000000c0200002100401000200000004000004200802000400000008000),
             .INIT_7A(320'h00000000021004010002000000000000000000000000000000108020080010000000000804200802),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000002100401000200000000200000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000210040100020000000000),
             .INIT_7D(320'h00000000000006200802000600000018000000000800000000000000040000400108020080010000),
             .INIT_7E(320'h00062008020006000062008020006000000000000000000000080200000000020000031004010003),
             .INIT_7F(320'h00062008020006000000000000000018802008001800000000180000000310040100030000000000)) 
           _a6640 ( .DOA({_d2961, _d2962, _d2963, _d2964, _d2965, _d2966, _d2967, _d2968, _d2969, _d2970, _d2971, _d2972, _d2973, _d2974,
                   _d2975, _d2976, _d2977, _d2978, _d2979, _d2980, _d2981, _d2982, _d2983, _d2984, _d2985, _d2986, _d2987, _d2988, _d2989,
                   _d2990, _d2991, _d2992, _d2993, _d2994, _d2995, na6640_36, na6640_37, na6640_38, na6640_39, na6640_40}),
                    .DOAX({_d2996, _d2997, _d2998, _d2999, _d3000, _d3001, _d3002, _d3003, _d3004, _d3005, _d3006, _d3007, _d3008, _d3009,
                   _d3010, _d3011, _d3012, _d3013, _d3014, _d3015, _d3016, _d3017, _d3018, _d3019, _d3020, _d3021, _d3022, _d3023, _d3024,
                   _d3025, _d3026, _d3027, _d3028, _d3029, _d3030, _d3031, _d3032, _d3033, _d3034, _d3035}),
                    .DOB({_d3036, _d3037, _d3038, _d3039, _d3040, _d3041, _d3042, _d3043, _d3044, _d3045, _d3046, _d3047, _d3048, _d3049,
                   _d3050, _d3051, _d3052, _d3053, _d3054, _d3055, _d3056, _d3057, _d3058, _d3059, _d3060, _d3061, _d3062, _d3063, _d3064,
                   _d3065, _d3066, _d3067, _d3068, _d3069, _d3070, _d3071, _d3072, _d3073, _d3074, _d3075}),
                    .DOBX({_d3076, _d3077, _d3078, _d3079, _d3080, _d3081, _d3082, _d3083, _d3084, _d3085, _d3086, _d3087, _d3088, _d3089,
                   _d3090, _d3091, _d3092, _d3093, _d3094, _d3095, _d3096, _d3097, _d3098, _d3099, _d3100, _d3101, _d3102, _d3103, _d3104,
                   _d3105, _d3106, _d3107, _d3108, _d3109, _d3110, _d3111, _d3112, _d3113, _d3114, _d3115}),
                    .ECC1B_ERRA({_d3116, _d3117, _d3118, _d3119}),
                    .ECC1B_ERRB({_d3120, _d3121, _d3122, _d3123}),
                    .ECC2B_ERRA({_d3124, _d3125, _d3126, _d3127}),
                    .ECC2B_ERRB({_d3128, _d3129, _d3130, _d3131}),
                    .FORW_CAS_WRAO(_d3132), .FORW_CAS_WRBO(_d3133), .FORW_CAS_BMAO(_d3134), .FORW_CAS_BMBO(_d3135), .FORW_CAS_RDAO(_d3136),
                    .FORW_CAS_RDBO(_d3137), .FORW_UADDRAO({_d3138, _d3139, _d3140, _d3141, _d3142, _d3143, _d3144, _d3145, _d3146, _d3147,
                   _d3148, _d3149, _d3150, _d3151, _d3152, _d3153}),
                    .FORW_LADDRAO({_d3154, _d3155, _d3156, _d3157, _d3158, _d3159, _d3160, _d3161, _d3162, _d3163, _d3164, _d3165, _d3166,
                   _d3167, _d3168, _d3169}),
                    .FORW_UADDRBO({_d3170, _d3171, _d3172, _d3173, _d3174, _d3175, _d3176, _d3177, _d3178, _d3179, _d3180, _d3181, _d3182,
                   _d3183, _d3184, _d3185}),
                    .FORW_LADDRBO({_d3186, _d3187, _d3188, _d3189, _d3190, _d3191, _d3192, _d3193, _d3194, _d3195, _d3196, _d3197, _d3198,
                   _d3199, _d3200, _d3201}),
                    .FORW_UA0CLKO(_d3202), .FORW_UA0ENO(_d3203), .FORW_UA0WEO(_d3204), .FORW_LA0CLKO(_d3205), .FORW_LA0ENO(_d3206),
                    .FORW_LA0WEO(_d3207), .FORW_UA1CLKO(_d3208), .FORW_UA1ENO(_d3209), .FORW_UA1WEO(_d3210), .FORW_LA1CLKO(_d3211),
                    .FORW_LA1ENO(_d3212), .FORW_LA1WEO(_d3213), .FORW_UB0CLKO(_d3214), .FORW_UB0ENO(_d3215), .FORW_UB0WEO(_d3216), .FORW_LB0CLKO(_d3217),
                    .FORW_LB0ENO(_d3218), .FORW_LB0WEO(_d3219), .FORW_UB1CLKO(_d3220), .FORW_UB1ENO(_d3221), .FORW_UB1WEO(_d3222), .FORW_LB1CLKO(_d3223),
                    .FORW_LB1ENO(_d3224), .FORW_LB1WEO(_d3225), .CLOCKA({_d3226, _d3227, _d3228, _d3229}),
                    .CLOCKB({_d3230, _d3231, _d3232, _d3233}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7378_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7379_10, na7380_9, na7382_10, na7383_9, na7384_10, na7386_9, na7387_10, na7388_9, na7390_10, na7391_9,
                   na7392_10, na7394_9, na7395_10, na7396_9, na7398_10, na7399_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7400_10, na7402_9, na7403_10, na7404_9, na7406_10,
                   na7407_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h6081014ba295810e8a528409014a106c992043a0e824294050e82528744695846908d214a1094202),
             .INIT_01(320'h15a52801a4e48049409694a0025a52801a42098210b920125025a006908260a029741d0745281082),
             .INIT_02(320'h841ac1304c1304c13050a48841304080a4d9741264ad2e8a50040842098210b920125020ad294004),
             .INIT_03(320'h84092e88501420480ba29745287452840842104c1405d0485480a508349014a106d2029420d24052),
             .INIT_04(320'h142049744280a1024ba2140508125d10a0284092e8850142049744280a1024ba2140508125d10a02),
             .INIT_05(320'h84210b4a500349c900928120214a1020ac00421085a52801a42001600210810841304080892e8850),
             .INIT_06(320'h300108421694a006939201250240429420494ba2300108421694a006939201250240429420415800),
             .INIT_07(320'h14a102104c1020220ac004210e48049409010a5081006042c0042106939201250240429420494ba2),
             .INIT_08(320'h812d294004b4a500348413042202149104c1405d14a52930509421d11a5611a4234090b485694a5d),
             .INIT_09(320'h910822108260850e02049439201250a4a0da4a5294a50641a4a5810b020d252922104c1085c90092),
             .INIT_0A(320'h9409680012870128125025a1005812834922401024a4694a5215a429085690a42208506c99204a54),
             .INIT_0B(320'h118128421c04a0494080b420604a0d2368495052210841305004042149b264a568581284a5d04052),
             .INIT_0C(320'h80a10210826084414a028105280a0414a0281202810841304080a5c95a52e82028364c802928125d),
             .INIT_0D(320'hb485210ad21484410a14b420084a4421044210842108413042812c0942502581284a04b025094096),
             .INIT_0E(320'h83204340c0900126c2c08320d21200812008125234a5290ad21484215a429084414a1024a4694a42),
             .INIT_0F(320'h810942104c1401004010040421745010210a41b480a5d040529420c843901420494086808126c2c0),
             .INIT_10(320'h143926c99214ba06021060210602106021060210602106021060210a4ba28419294ba2841b497450),
             .INIT_11(320'h6924483614803a0932529741214a5c90092812d280a5d1420d248906b04c1304c1304c1304c1304c),
             .INIT_12(320'h2104c1304c14050e824d8724024a14b4006102506925d0499294ba090a52e48049409694052e8a10),
             .INIT_13(320'h8745214852843a294a10e8a5087452843a29421d14a1d14a50e8a528108260a02e82c42098211010),
             .INIT_14(320'he8a429745297452e8a5d14ba297452e8a5d14ba29421d14a10e8a50874529421d14ac2843a290a50),
             .INIT_15(320'h83210e8a92e83a0e88841305014ba097412e825d04ba095204143a29421d04ba29585d1485290a10),
             .INIT_16(320'h60a02974528108260a029365d11a5611a42348528405d07412e825d04ba0974129741d04a1064190),
             .INIT_17(320'hb4a1625990b52029745285a42b0a16b42d215850b4a1690ad28589014a10258561420c8419081082),
             .INIT_18(320'h04ba2940842098280a9014a1024042b42d295850b020da40528409010ad0b4a56142c08349005a42),
             .INIT_19(320'he8a5080a10e82508744695846908d08108260a0294ba2940841305010b92b405d14a0225a5695a52),
             .INIT_1A(320'he8a5294a1d14a52943a294a0da13a097452843a294a10e825d07412e8a5d04ba297452843a097452),
             .INIT_1B(320'h2098280a4d932560321d04ba08744695846908d0e48149409605a029745d04ba294a528745294a50),
             .INIT_1C(320'h14a10e8252e8a5d14a10e8252e8a508741297452843a094ba29421d04a5d14a10e8252e83a294204),
             .INIT_1D(320'h04a5297452843a094a52e8a508741294a5d14a10e8252e8a5d14a10e8252e8a5d14a10e8252e8a5d),
             .INIT_1E(320'h10a5081040b00108409010a50810560021084a528124413042240429420405800842149104c1405d),
             .INIT_1F(320'h14a50e8892e8a502104c1405d058841304220204209826098280ba094a50e825294a042104c10890),
             .INIT_20(320'h14a10e8a52843a2958508745214a10e8a4290a50874529421d14a10e8a5087452843a2943a294a1d),
             .INIT_21(320'h94ba297452e8a5d14ba297452e8a5d14ba297452e8a5d14ba297452e8a5d14ba297452843a29421d),
             .INIT_22(320'h34ac2348468409034ac2e8a50e825d04ba097412e825d14a10e825d14ac2e8a42948508745214ba2),
             .INIT_23(320'h04ba097412e825d04a5d0741284192040842108413050148901745287456e8ad2b0ad215a90243a2),
             .INIT_24(320'hb1a10042008348484852b5ad234856840108020c840102405d14a0d9744695846908d214a101741d),
             .INIT_25(320'h14a10e8192043a234ac2348468408414a04852029420cb324264850040900408484852b5ad234856),
             .INIT_26(320'he8242843a090a1690ad2843a0974042098280a5d14a04209828020080a4d9744695846908d081202),
             .INIT_27(320'h8405285a508021094a160021087412240429421d04a1680a10e8242843a094ba090a10e8242843a0),
             .INIT_28(320'h80a5d102c0812d011a02b4a0297440b0214910522108260a0297412e88d2b08d211a4294a1694200),
             .INIT_29(320'h210842129220a442098280ba297452e8a5d14ba297452e8a4420982112441304080896808d015a52),
             .INIT_2A(320'he8a5d14ba297452e8a5d1489295a0214a52b0a0d24a568085614192012c0b400497444974449744d),
             .INIT_2B(320'he8a5d14a16e8a5d14ba2942dd14ba297452858869364cb4056143a29349491084130501438081250),
             .INIT_2C(320'h14052974528108260a021725680ba294044b4ad2b4a4097452810841305017452e0204943a297452),
             .INIT_2D(320'h8741297452e8a508741297452843a094ba29421d04a5d14a10e8252e8a50874129741d14a102104c),
             .INIT_2E(320'h94ba29421d04a5297452843a094a52e8a508741297452e8a508741297452e8a508741297452e8a50),
             .INIT_2F(320'h8408205800842048085284082b00108425294092209821120214a10202c004210a488260a02e8252),
             .INIT_30(320'h1125d14a042108260a02e82c420982110102104c1304c1405d04a528741294a50210826084480852),
             .INIT_31(320'h14a5087452b0a10e8a429421d1485214a10e8a52843a29421d14a10e8a508745287452943a294a1d),
             .INIT_32(320'he825d04ba097412e8a4297452843a097452b0ba290a521421d14852e8a52e8a5087452843a29421d),
             .INIT_33(320'h14052e8a502104c14052e8ad2b0ad215ba02104c140101488484852e8a50e8ad2b0ad215ba097412),
             .INIT_34(320'h832526484c90a00840102121214ba2943a0958c424242974528744695846908d024ba0210842104c),
             .INIT_35(320'h802100408484ad6308d214ad6308d2b58c23401080210041a42424295ac611a56b18468021004200),
             .INIT_36(320'h95a5204ba294084209828020080a5c900928744695846908d0b020d274569585690ad21108424010),
             .INIT_37(320'he8252e8a508741297452843a094ba0e8a508108260a0294ba2940841305010b92b405d14a0225a56),
             .INIT_38(320'h94ba297452843a094ba297452843a094ba297452843a094ba297452843a094ba29421d04a5d14a10),
             .INIT_39(320'h9104c1089010a50810160021085244130501741294a5d14a10e825294ba29421d04a5297452843a0),
             .INIT_3A(320'h2108260a02e8252943a094a5281084130422404294204102c0042102404294204158008421294a04),
             .INIT_3B(320'h943a294a1d14a042098280ba234ac23484614a0085204942928745210250e8a5294050e8a5294050),
             .INIT_3C(320'h9409680252e8a50693a087452943a2940842104c14050e8a5025a0294ba29409680a52e8a5024ba2),
             .INIT_3D(320'h2108420880912c413084130106c98660192b3046e4812670422304ce48422418260a02e8a50e4004),
             .INIT_3E(320'h9108421084210841304080204833a420a42b4acc919922125624ba4210842085210a442104c143a4),
             .INIT_3F(320'h240842108421084210826080280200802100439c65042119829485d908429764290a521498290852),
             .INIT_40(320'hb08c260992931a2689a21379280990b499293252148429084290852b364ce0a0c941926004293240),
             .INIT_41(320'h1324de4b8d3198260a5295a5264992948521084c6498c631a26498d908cd1484c60a12634461184d),
             .INIT_42(320'h80202e7040859a2688c6e099c141b29745264a52b30506c89294190b4a5664a526ca4d13442649a2),
             .INIT_43(320'h94842134426884c9724093652036dd14a4c9304c91a5211ad6b325004a4c9324c100500401004010),
             .INIT_44(320'h1084c1725c90a526884d1325c9024d9480d949a21439c141b2e4a4c936521365294996940129324c),
             .INIT_45(320'he085069a463324cb584ce7050608c6e4810e7084141bc93642b199264992134426898c1084260982),
             .INIT_46(320'hb4acc919922125624bb22104290852210826f2dce08506f38085a526f382141a28098213052e49bc),
             .INIT_47(320'h97444209828779d20982040102199d2105215a5624ac497482148521108413050040102419d20a42),
             .INIT_48(320'h30b9614ad23184614852b18c293182b7452e884c130842104c1400687452ec8442104c10050e8a4c),
             .INIT_49(320'h1744cb0ac214ac290992609969488421084b584221a421198201a06e98843585630a4d1304080050),
             .INIT_4A(320'h040d66344c348c294842b5ac6b0a4c3585d132cc15996b18c61304cb58d6b4a46b1ac21744c11ac2),
             .INIT_4B(320'h948843488421046348961488269b9c6f38d059a2171a637242b4a4c959b268986634c66305004010),
             .INIT_4C(320'h318423185d1325231842e898294b9c69b8c682dc331a6332cc1020080200140d661ad2b324c34a46),
             .INIT_4D(320'h2125634896148826885c69a421344261ac6b5ad635a5c9184c6c8d2149a26d982932d210add91a46),
             .INIT_4E(320'h64a463085d13052934cc6f19c682dc331a6332cc1020080200140d6658d2b324cb48469488434884),
             .INIT_4F(320'h10982b7642908c297646903a490a4614bb23485d90a4230a5d91a42e9a42148d690ac6b585630ba2),
             .INIT_50(320'h2184694add10a52e8a42210842124214884b58841188269ad6b0a42171a6e88521344d35992948dd),
             .INIT_51(320'h00a0217452213b26319290844210842108260a16802008020000a50e8a56b7452b4bb2308d2b4a1d),
             .INIT_52(320'h3498d318c6b184213484e3246e8a5d134dd11096630d268a4427452631cc609a22118c1024080210),
             .INIT_53(320'h10856b58c691a46358d63485231842948423185635acc9305211ba297442698c6b5a5d172442598c),
             .INIT_54(320'h308c080ad634982b4ba2b199211084131a42344214b8210b9237452e89a6b58c615a4d3185213386),
             .INIT_55(320'h93252609b2971b2618c2b1ad6930461184085ac693056974442098c13652e364c3185635ad260a06),
             .INIT_56(320'h35a52b5986130d6930d234acc1498c10a4214992931a693050e9ad26184430846609869304c10a52),
             .INIT_57(320'h109a2618c6b1a421485610856b0842b584215a52949863098610ac610842b58c294a46b184211856),
             .INIT_58(320'h6419090a46b1ac0b1056690962420c94a1c80842b08c6302cc60992902cd948cc1318293050043a4),
             .INIT_59(320'h031c42184660046601c27700c309d2942cc31810b199c1018404a4611b8061a02b39a494a0485a0c),
             .INIT_5A(320'h912d2959ce60850e904234992670168598e9798283a5ee905215992b1056202c4b12c4b12cd2599c),
             .INIT_5B(320'heca42340dd21042337a275a56734d2e32169325d130408020083246908d677884210841364c731cc),
             .INIT_5C(320'h1c0d68ca74b59b2b34423401d9484685b92808c4b0b92808c4b088694a4c1481620add108d2b3250),
             .INIT_5D(320'hf7bdef7bdef7bdefffdef7bdef7bdef7bdefffdef7bdef7bdef7bdefffdef7bdef7bdef7bde0782b),
             .INIT_5E(320'hf7bdef7bdef7bdefffdef7bdef7bdef7bdefffdef7bdef7bdef7bdefffdef7bdef7bdef7bdefffde),
             .INIT_5F(320'h294a55000000000500000000057bdef7bde518c6318c655ad6b5ad6fffdef7bdef7bdef7bdefffde),
             .INIT_60(320'h6318d711ca635cd721ed6b5406b88e4812e694ac03529500000000050000000005000000000514a5),
             .INIT_61(320'h6b1cc7118d431cd6b1cc639aa235a42388d735446918c731ac700ee6380d638ae635ae23944611c4),
             .INIT_62(320'h5192d7394e231ac6a809734c52b00e719ad739ca00000061ef7bcc353c3c8208d6908e2118d431cd),
             .INIT_63(320'h2214848000635cc6288d7218a5012c739ce700ce7380a718c52b00d5910a42408021ac6110d6308e),
             .INIT_64(320'h210810916c205cc031800000000000500a6295806ac8852120221092288a211083280a618a5601ab),
             .INIT_65(320'h435cc6a9c46398d531cc731aa02986314ac6a1cc711ca080046908b029cc2958f63084691ad030ec),
             .INIT_66(320'h631ce235cd6b98e500c43b1cd231a83b484539847b58e6b98c6908a235c8231c8090c77390c6b88e),
             .INIT_67(320'h33ade0a639022189ec6b9684aaf4ada708cfdde7f59c6cc521c4100025ed6b18d7200a7318c614ac),
             .INIT_68(320'hbfcef860088e42912a5a1ae7b2329c2b6bd71bd679ff7403104873158f7350b52697b5613943beff),
             .INIT_69(320'h0000000000000000000000000331a4235004b9ed694ac735ce735ced4942dcd63e5184ed5a5b78ce),
             .INIT_6A(320'h6390c5314891801025cd721cc295806bdce6b9af7395194e96b00210842108421084200000000000),
             .INIT_6B(320'h4ad447110042d447110042d44711014a96a238885318d238880388c6a8880398a4a02e638887054c),
             .INIT_6C(320'hb01b80018d7118a221895112a0b1ac69d00711cc3a084731ce4b1a46b9c42200e639074058d628e8),
             .INIT_6D(320'hf7bfff7bdef7bdef7bdef7b57400013b00a680ee22809739af734a56380721dcc6b9ae403c158e06),
             .INIT_6E(320'hf7bfff7bdef7bdef7bdef7bfff7bdef7bdef7bdef7bfff7bdef7bdef7bdef7bfff7bdef7bdef7bde),
             .INIT_6F(320'hb5bfff7bdef7bdef7bdef7bfff7bdef7bdef7bdef7bfff7bdef7bdef7bdef7bfff7bdef7bdef7bde),
             .INIT_70(320'h0014000000001400000000145294a5295400000000140000000015ef7bdef7946318c631956b5ad6),
             .INIT_71(320'h7908e525c86a9ac239aa0118d735cc631a6700e43b98d735c8711ce0258c630a5601a12294000000),
             .INIT_72(320'h868000398e0108743d4d435c42318c7280a6848d43984531004b9cd7b0c52b00d711ce6bf000014d),
             .INIT_73(320'haef7bd6f78080c6731ae611c902d046a48e4818d211c90b88e4818a620ac739cc610246a585034ba),
             .INIT_74(320'h00000000000000000000000000000000000067a000000ea5c949e294a5293252949975def3bbef7b),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6641 ( .DOA({_d3234, _d3235, _d3236, _d3237, _d3238, _d3239, _d3240, _d3241, _d3242, _d3243, _d3244, _d3245, _d3246, _d3247,
                   _d3248, _d3249, _d3250, _d3251, _d3252, _d3253, _d3254, _d3255, _d3256, _d3257, _d3258, _d3259, _d3260, _d3261, _d3262,
                   _d3263, _d3264, _d3265, _d3266, _d3267, _d3268, na6641_36, na6641_37, na6641_38, na6641_39, na6641_40}),
                    .DOAX({_d3269, _d3270, _d3271, _d3272, _d3273, _d3274, _d3275, _d3276, _d3277, _d3278, _d3279, _d3280, _d3281, _d3282,
                   _d3283, _d3284, _d3285, _d3286, _d3287, _d3288, _d3289, _d3290, _d3291, _d3292, _d3293, _d3294, _d3295, _d3296, _d3297,
                   _d3298, _d3299, _d3300, _d3301, _d3302, _d3303, _d3304, _d3305, _d3306, _d3307, _d3308}),
                    .DOB({_d3309, _d3310, _d3311, _d3312, _d3313, _d3314, _d3315, _d3316, _d3317, _d3318, _d3319, _d3320, _d3321, _d3322,
                   _d3323, _d3324, _d3325, _d3326, _d3327, _d3328, _d3329, _d3330, _d3331, _d3332, _d3333, _d3334, _d3335, _d3336, _d3337,
                   _d3338, _d3339, _d3340, _d3341, _d3342, _d3343, _d3344, _d3345, _d3346, _d3347, _d3348}),
                    .DOBX({_d3349, _d3350, _d3351, _d3352, _d3353, _d3354, _d3355, _d3356, _d3357, _d3358, _d3359, _d3360, _d3361, _d3362,
                   _d3363, _d3364, _d3365, _d3366, _d3367, _d3368, _d3369, _d3370, _d3371, _d3372, _d3373, _d3374, _d3375, _d3376, _d3377,
                   _d3378, _d3379, _d3380, _d3381, _d3382, _d3383, _d3384, _d3385, _d3386, _d3387, _d3388}),
                    .ECC1B_ERRA({_d3389, _d3390, _d3391, _d3392}),
                    .ECC1B_ERRB({_d3393, _d3394, _d3395, _d3396}),
                    .ECC2B_ERRA({_d3397, _d3398, _d3399, _d3400}),
                    .ECC2B_ERRB({_d3401, _d3402, _d3403, _d3404}),
                    .FORW_CAS_WRAO(_d3405), .FORW_CAS_WRBO(_d3406), .FORW_CAS_BMAO(_d3407), .FORW_CAS_BMBO(_d3408), .FORW_CAS_RDAO(_d3409),
                    .FORW_CAS_RDBO(_d3410), .FORW_UADDRAO({_d3411, _d3412, _d3413, _d3414, _d3415, _d3416, _d3417, _d3418, _d3419, _d3420,
                   _d3421, _d3422, _d3423, _d3424, _d3425, _d3426}),
                    .FORW_LADDRAO({_d3427, _d3428, _d3429, _d3430, _d3431, _d3432, _d3433, _d3434, _d3435, _d3436, _d3437, _d3438, _d3439,
                   _d3440, _d3441, _d3442}),
                    .FORW_UADDRBO({_d3443, _d3444, _d3445, _d3446, _d3447, _d3448, _d3449, _d3450, _d3451, _d3452, _d3453, _d3454, _d3455,
                   _d3456, _d3457, _d3458}),
                    .FORW_LADDRBO({_d3459, _d3460, _d3461, _d3462, _d3463, _d3464, _d3465, _d3466, _d3467, _d3468, _d3469, _d3470, _d3471,
                   _d3472, _d3473, _d3474}),
                    .FORW_UA0CLKO(_d3475), .FORW_UA0ENO(_d3476), .FORW_UA0WEO(_d3477), .FORW_LA0CLKO(_d3478), .FORW_LA0ENO(_d3479),
                    .FORW_LA0WEO(_d3480), .FORW_UA1CLKO(_d3481), .FORW_UA1ENO(_d3482), .FORW_UA1WEO(_d3483), .FORW_LA1CLKO(_d3484),
                    .FORW_LA1ENO(_d3485), .FORW_LA1WEO(_d3486), .FORW_UB0CLKO(_d3487), .FORW_UB0ENO(_d3488), .FORW_UB0WEO(_d3489), .FORW_LB0CLKO(_d3490),
                    .FORW_LB0ENO(_d3491), .FORW_LB0WEO(_d3492), .FORW_UB1CLKO(_d3493), .FORW_UB1ENO(_d3494), .FORW_UB1WEO(_d3495), .FORW_LB1CLKO(_d3496),
                    .FORW_LB1ENO(_d3497), .FORW_LB1WEO(_d3498), .CLOCKA({_d3499, _d3500, _d3501, _d3502}),
                    .CLOCKB({_d3503, _d3504, _d3505, _d3506}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7415_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7416_10, na7418_9, na7419_10, na7420_9, na7422_10, na7423_9, na7424_10, na7426_9, na7427_10, na7428_9,
                   na7430_10, na7431_9, na7432_10, na7434_9, na7435_10, na7436_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7438_10, na7439_9, na7440_10, na7442_9, na7443_10,
                   na7444_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h0048029c0529ce7014a739ca7b9ce701ec739c05014a639ce7014a73c0b52d4d631ee7420e731ce7),
             .INIT_01(320'h39ee739c0cf1cee39c87b9ce721ee739c0e30401003c73b8e719ce7038c100405380a0280a7399c1),
             .INIT_02(320'h39c023a0e43b0ec388e729cce08024014e0380a565ee7014e721ccc70401003473b0e701cf739ce4),
             .INIT_03(320'h39c078148739ce039e05380a7380a739c866382008000294043dce738087b9ce700cf739ce019ee7),
             .INIT_04(320'h39ce0380a439ce701c0521ce7380f0290e739c078148739ce03c0a439ce701e0521ce7380f0290e7),
             .INIT_05(320'h39ce63dce73809c39cc73c8f7b9ee705cf739ce731ee739c0601ce7b9ce73998e080240000701487),
             .INIT_06(320'h25ce739cc7b9ce7002c7388e791ef73dce0b9c0525ce739cc7b9ce700b87390e791ef73dce0b9ee7),
             .INIT_07(320'h294e7318200900001cf739ce791cee39e47bdcf7380e7398f739ce703ac7380e791ef73dce0b9c05),
             .INIT_08(320'h390f739ce43dce7381c60802039ce53982008000296f73d0e731ce02d4b5358c7b9dd73dcf735ce0),
             .INIT_09(320'h331c4110c1004a761cec39f473a8e77dce07dee7bdee7a1c0a79ce739ce063c67218200801e39dc7),
             .INIT_0A(320'h39c0731ce7388e7398e701ce639ce7380c701ce711ce1bdce7b9ef618f08c59ce218c601cc6310cb),
             .INIT_0B(320'h290e7398e239cec39c07398e739ce0601e338ce721886080242002509c0735ee739ce7398f0294d7),
             .INIT_0C(320'h39ce7710c100400b9cf7382e73dce0b9cf7380f73888608024014f6bdce7814a6380e639de7380e0),
             .INIT_0D(320'h1ceca579deb2d62318c5318c6310c22188e008864298e080253b8e7b9ce771cf739cee39ee739dc7),
             .INIT_0E(320'h3b0e0398e731ce701ce73b0e0300e7380e73b0e70dee73dcf7b3de6c23164a4ce318c6018c1b58d3),
             .INIT_0F(320'h3f987338200ad6a5252420020080a531ce701c0039cf0294d739cec39d0739ce639c0731ce701ce7),
             .INIT_10(320'h39e4701cc739e0511ce751ce711ce751ce711ce751ce711ce751ce739c0539dd739c0539c07380a7),
             .INIT_11(320'h008ec380ec39e052a2f73c0a5318f239c87390e739cf029ce021d87008e8398e03b8e8398ee3b8e8),
             .INIT_12(320'h2182000000080a7014a03d0e701cec398e739ce7000f029517b9e05298c791ce239c8739ce7814e7),
             .INIT_13(320'h3c0a5318e739e0529ce7814e73c0a739e0539cf029cf0294e7814a7399c100400816a670401000e7),
             .INIT_14(320'h014a6380a53c0a5814b0296052c0a5814b02960529cf0294e7814a73c0a539cf0296e739e05298e7),
             .INIT_15(320'h3e0e7815e701405814c60802029c05280a5014a029405284e139e0529ce0294052dce0294c731ce7),
             .INIT_16(320'h004053c0a7399c100405380f02d4b5358c7b9d08b9ce0280a5014a029405280a5380a0296e741cc7),
             .INIT_17(320'hb98e741d87384f73c0a5b9ee7b98e735cf73dcc739ae7b9ee639c27b9ce701ee739ce439e07399c1),
             .INIT_18(320'h39a0539c863040100027b9ce781ef73dcf735cc73dce009ee739e07bdcf73dcd731cf738207b9ee7),
             .INIT_19(320'h814b739ce7014b73c0b52d4d631ef7398c10040539e0539cce0802000217b9cf029ce071ee7b9ee7),
             .INIT_1A(320'h814b7bdcf0296f7b9e052dce06ba05280a539c0529ce7814a02c0a5814b0296052c0a739e052c0a5),
             .INIT_1B(320'h70401014e03d8e73a8e0294052c0b52d4d631ee7e1ced39dc73dcf73c0b0296052def73c0a5bdee7),
             .INIT_1C(320'h29ce7014a7814f029ce7014a7814e7380a53c0a739c0529e0539ce0294f029ce7014a78160539ce6),
             .INIT_1D(320'h296f73c0a739c052dee7814e7380a5bdcf029ce7014a7814e029ce7014a7814f029ce7014a7814f0),
             .INIT_1E(320'hbdcf7382f73dce739e47bdcf7382e7b9ce73dad7bd4e60802091ef73dce039ee739ce53982008000),
             .INIT_1F(320'h294e7814c7014e733820080102d4ce0802001ce43040000001002052dee7814b7bdce43382008247),
             .INIT_20(320'h294e7014a739c052dce73c0a531ce7814a631ce73c0a539ce029ce7014e7380a739c0539c0529ce0),
             .INIT_21(320'h29e052c0a5814b0296052c0a5814b0296052c0a5814b0296052c0a5814b029605280a539c0529ce0),
             .INIT_22(320'ha96a6b18f7b9c4739ee7014e7014a029405280a5014a0294e7014a0294e7014a6398e73c0a531e05),
             .INIT_23(320'h29405280a5014a0294e0280a5b9f0739cce008860802029cc7380a73c0b7816e5b9ae63dd27c1e05),
             .INIT_24(320'h318c6318e7381cc31ce639aa532526318c639cee39ce741ce029ce03c0b52d4d631ee7422e7380a0),
             .INIT_25(320'hb9ee701407b9c05a96a6b18f739dcc398f83a4f739ce4be0c6618c739cc739dcc31ce639aa531086),
             .INIT_26(320'h014a6b9c05298e7b9ee6b9c05280a670401014e029ce6704014a484014e0380b52d4d631ef73e0f7),
             .INIT_27(320'h39cd739cf739ce735ce7b9ce7380a5c1ef73dce0294e739ee7014a6b9c0529c0529ae7014a6b9c05),
             .INIT_28(320'h3dce0290e7b80e6b9ef7bdcf7380a439ee43d4e7331c100405380a5016a5a9ac63dce845ce73dce7),
             .INIT_29(320'h25d8e00887a9ce67040100005280a5014a029405280a5014a670401054e6080240000735cf7bdcf7),
             .INIT_2A(320'h014a029405280a5014a0296f7bdef7b9ef7b9ce0bdee7bdef739f073b0e739cee380a0380a2380a0),
             .INIT_2B(320'h014a0294e7014a02940529ce029405280a539c47380e6b9cf739c05281c3390c6080202dd07390e7),
             .INIT_2C(320'h080a73c0a7399c100400042f739e0539c0e3dcf73dce7340a7390c608020000a501cee39c05280a5),
             .INIT_2D(320'h380a5380a7014e7380a5380a739c0529c0539ce0294e029ce7014a7014e7380a53c0a029ce733820),
             .INIT_2E(320'hb9c0539ce0296f7380a739c052dee7014e7380a5380a7014e7380a5380a7014e7380a5380a7014e7),
             .INIT_2F(320'hb9c17b9ee739cf03dee7b9c173dce739ed6bdea730401040f7b9ee701cf739ce729cc100400014b7),
             .INIT_30(320'h298f029ce6531c100400816a670401000e7218200000008010296f73c0a5bdee7219c1004103dee7),
             .INIT_31(320'h294e73c0a5b9ce7014a639ce0294c639ce7814a739e0539cf029ce7814e73c0a73c0a539e0529cf0),
             .INIT_32(320'h014a029405280a5014a63c0a539c052c0a5b9e05298e639ce0294c7014a7814a73c0a539e0529cf0),
             .INIT_33(320'h080a7814e733820080a7016e5b9ae63dc05338200908029dcc39087814e7016e5b9ae63dc05280a5),
             .INIT_34(320'h3a0e6c14a4294e7398c7100e421e0539c0529cce61d293c0a7380b52d4d631ee721c057380221820),
             .INIT_35(320'h39ce529d4831cc7c20e5298e6c20c5316632a105318c739c0a418e731cd8418a62cc65420a6318e7),
             .INIT_36(320'hb9ee739a0539c86304014a484014fa3dee7bc0b52d4d631ee739ee0bc0b72dcd731ee840806218c6),
             .INIT_37(320'h014a7814e7380a53c0a739c0529e05814e7399c10040539e0539cce0802000217b9cf029ce071ee7),
             .INIT_38(320'h29e05380a739c0529e05380a739c0529e05380a739c0529e05380a739c0529c0539ce0294e029ce7),
             .INIT_39(320'h3982008387bdcf7380e7b9ce7394e608020000a5bdcf029ce7014b7b9e0539ce0296f73c0a739c05),
             .INIT_3A(320'h218c100400814b7b9e052def7390ce08020e1ef73dce0bdcf739ce7e1ef73dce0b9ee739cf6b5ef5),
             .INIT_3B(320'h39c0529ce029ce63040100205a96a6b18f7420c73b8efb9df7380a5b9ce7014b7b9ce7014b7b9ce7),
             .INIT_3C(320'h39da739cc7014e703a05280a539c0539c4431820080a7014e771ce7b9c0539dc739ee7014e771c05),
             .INIT_3D(320'h731067188528aea080083a0e781c05b1cc7280a5e1ce70686602860b146600dc300400014e711cee),
             .INIT_3E(320'hb8886510c863802080292100039800614a621cf439d87510e719e06201c6114c5490801102008006),
             .INIT_3F(320'h11dc0110ca6380221901005256316b529242025433c89a12ca4ad90314d42c0a53199a5d0cb22549),
             .INIT_40(320'h6dcf765d973a204812042034b490073dc973a0cf7b9c3420a62914db40a8024be5a70b61589212eb),
             .INIT_41(320'h212f001c80526441512c2668491ec6b9ceda529a01c8c61a04e5f50211505108ae1cf2e408ab9ef0),
             .INIT_42(320'h21009a008529e048292a311c029604640a5216e9cd9a98258461c0739af641ae7834902408425e04),
             .INIT_43(320'hb9a94a42b5856a8b9985bc2ac280903188e21a9ad1f57214a5bf1852d086b8ae00a4ad6b18b5a949),
             .INIT_44(320'hef7a0bd88ad5357856b0a9ae6616f02b0b049a05495c029606018fc3c1262409ad5cc7614b421ae2),
             .INIT_45(320'h015250288a4f1243b538500a57112471ce71008629608b80e46930d65e97241a401386bf7bdc1384),
             .INIT_46(320'h21cf439d87510e719e09718a62a48442981810e8024a58600529ce984809296092949d2d0b775e14),
             .INIT_47(320'h3c08620401041d03040149080010d0628a531ce721ce33c0c53152420044080294908001cd0614a6),
             .INIT_48(320'h25f46a1ed621ee6b5885b5ce73b187380a4024a0208022182009085000a50108221820090a0814b8),
             .INIT_49(320'h280bea6b34b9094524ca621862a0443298e2dd25458e70a00121405810c4294252def020029210a0),
             .INIT_4A(320'h200a5c00bc29c94a52e4252e7b9ce2250a02f8ec29347bdee7390e232b474df2a31e87280be39324),
             .INIT_4B(320'h3988ea6402331292d1073d1418574c840d02de152c2052f0e4252fab920781549d40a5c002a52524),
             .INIT_4C(320'h29b2aca8a02faf756d45017cabdd4c81118812fc272042e2e00ad4a4a48428087e1ac73d0c6ce55b),
             .INIT_4D(320'h010842e4473e5c1854b281ef7bc085914f7358b6ad4e4298c6858e7bd60a81ec63c0e63d8e0294c6),
             .INIT_4E(320'hf5eeaca8a02f957bc09681ac4812fc272042e2e00ad4a4a48428087e1ac73d8c6a697939986a690a),
             .INIT_4F(320'hc978a380a5358b5a80a531806294c6b5405298c0294c656aa0294c6024a531949d193621d5451405),
             .INIT_50(320'h310b4adc80290bc06d4950048638a552486dd1ca63181810944d73ad6205064a5d415021f474a4a0),
             .INIT_51(320'h21409240a51020557b4952880429c221981004856316b52929214a0014a4200bb21414216975f0a0),
             .INIT_52(320'hb9f402ee95b94a63c040568e7014802c2802881744ae7814a0140a565014e2604100c00a4ab52924),
             .INIT_53(320'h2d0e6ad8d6b12c4b1c8645ed62aebbad8882ecd6adcca3a0c6394052016586494b9ce02b8e205d10),
             .INIT_54(320'h2d4a401ce7a1dc739c05212c4218440aa02040e559e4629d87380a4016153de9629cf0492f7ccb4b),
             .INIT_55(320'h290a6016173ea07b1e8739ee738025a94e401cf43a8e738086205402c2e7b40f63d0e73dce700485),
             .INIT_56(320'h39cf6b1815382a73a8a7a9caa29c02298b7b9e873021538020054e7014e6a84e8017453f0e429af7),
             .INIT_57(320'h38607014f5396e5b1ed7bdee6bdef735ef7bded6b580539485b5ae6b96f735cc6b5ac7b98d7bdcf7),
             .INIT_58(320'h21cc7298c7a9ac53a0f780008521ccb9cf43b90529915b0ce095f1731ed0bd4a4b8285380252820e),
             .INIT_59(320'h3020601ce731cf7d1e18338c63d8d7398a0a94a739c1c29c082dce739dc7318f731e04b9ce039ce0),
             .INIT_5A(320'hb80e7b1e07004a0018a1a96c7078e639c1039c01040e7018a5095473a8f741ee4398e83a8f005c1e),
             .INIT_5B(320'h056a5a9680218a1ac00585cf73c287028e7b88b02802a4a4840489a4a68421c864298e0c0a080006),
             .INIT_5C(320'h00c0418c6319205a8025a8080ad4b52dd9739ee4b9d9739ee4b9d17bdcf4b9cf701ee029aa5acae7),
             .INIT_5D(320'h294a5294a5294a5084a5294a5294a5294a5084a5294a5294a5294a5084a5294a5294a5294a500402),
             .INIT_5E(320'h294a5294a5294a5084a5294a5294a5294a5084a5294a5294a5294a5084a5294a5294a5294a5084a5),
             .INIT_5F(320'h0000008000000000842108421080000000008000000000800000000084a5294a5294a5294a5084a5),
             .INIT_60(320'h992602dd34224144e0a1748a0d2529281c07366f0040108000000000800000000084210842108000),
             .INIT_61(320'ha326441a4ea8105a32646bdd229c17294217ba45294bf9035f90009fc8007200090005ba684a3124),
             .INIT_62(320'ha006e28288349897140e81e099bc019006e0c8b400000014842124e51126294a705ca50ca4ea8105),
             .INIT_63(320'h811eb780102b0a0d0494a10ef281c0086d428313a140103a049bc0e0408f5bc0103cee2a5e771529),
             .INIT_64(320'h4a52a2a6cf27489018c000000000000807984de0702047ade0c0093c030009816bb40184693781c0),
             .INIT_65(320'h4d006714a5a00ce2cc03295c5016159366f030b34193449433acca50061924df52e486711af00000),
             .INIT_66(320'h748b424c05a2705a0318000139500c414c82801500188c9860999050500604c0600300094b43d468),
             .INIT_67(320'hd6b5a4a52942108bdef7b5ad6294a5210849ce7394a520842100000038a1716744e001849ce9166f),
             .INIT_68(320'h5ad6bc6318ce739318c639ce7a5294ad6b51084218c63842108c631ffffff7bde6b5ad6318cdef7b),
             .INIT_69(320'h0620800018862080201882000c1002401807428e9366f049a5049a5739ce7bdefe739cef7bd5294a),
             .INIT_6A(320'h73dce29de20902103a144e25694de070428701b04b52318c63200188620802018820000621882008),
             .INIT_6B(320'h914290b440f90290b440f90290b4404fe81485a2a00a0305a201603002a2015d5288059d262a80b4),
             .INIT_6C(320'h20715000ac2b0ef24984292a905093914404d13200aac2bc3a0029029534688054824e101ee75002),
             .INIT_6D(320'h29421294a5294a5294a5296d59800028405080a1b140e039b07a6b37d4059152448289c002010060),
             .INIT_6E(320'h29421294a5294a5294a529421294a5294a5294a529421294a5294a5294a529421294a5294a5294a5),
             .INIT_6F(320'h00021294a5294a5294a529421294a5294a5294a529421294a5294a5294a529421294a5294a5294a5),
             .INIT_70(320'h00020000000002108421084200000000020000000002108421084200000000020000000002000000),
             .INIT_71(320'h560a71cea0a16ba195d503255ab82e9cdd0a80b22a48905138a4d3503a0e91533781c02a42000000),
             .INIT_72(320'h9c00001432060a0200206540566a80a5005080a0655432baa0701cd84e099bc0ea4d3530fe0000a1),
             .INIT_73(320'h00000000000029a29dc148e5904565184b2c834f90e5903932c8041025408ce401114493a86025d3),
             .INIT_74(320'h0000000000000000000000000000000000001ce0000001904421084210841908420c400000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6642 ( .DOA({_d3507, _d3508, _d3509, _d3510, _d3511, _d3512, _d3513, _d3514, _d3515, _d3516, _d3517, _d3518, _d3519, _d3520,
                   _d3521, _d3522, _d3523, _d3524, _d3525, _d3526, _d3527, _d3528, _d3529, _d3530, _d3531, _d3532, _d3533, _d3534, _d3535,
                   _d3536, _d3537, _d3538, _d3539, _d3540, _d3541, na6642_36, na6642_37, na6642_38, na6642_39, na6642_40}),
                    .DOAX({_d3542, _d3543, _d3544, _d3545, _d3546, _d3547, _d3548, _d3549, _d3550, _d3551, _d3552, _d3553, _d3554, _d3555,
                   _d3556, _d3557, _d3558, _d3559, _d3560, _d3561, _d3562, _d3563, _d3564, _d3565, _d3566, _d3567, _d3568, _d3569, _d3570,
                   _d3571, _d3572, _d3573, _d3574, _d3575, _d3576, _d3577, _d3578, _d3579, _d3580, _d3581}),
                    .DOB({_d3582, _d3583, _d3584, _d3585, _d3586, _d3587, _d3588, _d3589, _d3590, _d3591, _d3592, _d3593, _d3594, _d3595,
                   _d3596, _d3597, _d3598, _d3599, _d3600, _d3601, _d3602, _d3603, _d3604, _d3605, _d3606, _d3607, _d3608, _d3609, _d3610,
                   _d3611, _d3612, _d3613, _d3614, _d3615, _d3616, _d3617, _d3618, _d3619, _d3620, _d3621}),
                    .DOBX({_d3622, _d3623, _d3624, _d3625, _d3626, _d3627, _d3628, _d3629, _d3630, _d3631, _d3632, _d3633, _d3634, _d3635,
                   _d3636, _d3637, _d3638, _d3639, _d3640, _d3641, _d3642, _d3643, _d3644, _d3645, _d3646, _d3647, _d3648, _d3649, _d3650,
                   _d3651, _d3652, _d3653, _d3654, _d3655, _d3656, _d3657, _d3658, _d3659, _d3660, _d3661}),
                    .ECC1B_ERRA({_d3662, _d3663, _d3664, _d3665}),
                    .ECC1B_ERRB({_d3666, _d3667, _d3668, _d3669}),
                    .ECC2B_ERRA({_d3670, _d3671, _d3672, _d3673}),
                    .ECC2B_ERRB({_d3674, _d3675, _d3676, _d3677}),
                    .FORW_CAS_WRAO(_d3678), .FORW_CAS_WRBO(_d3679), .FORW_CAS_BMAO(_d3680), .FORW_CAS_BMBO(_d3681), .FORW_CAS_RDAO(_d3682),
                    .FORW_CAS_RDBO(_d3683), .FORW_UADDRAO({_d3684, _d3685, _d3686, _d3687, _d3688, _d3689, _d3690, _d3691, _d3692, _d3693,
                   _d3694, _d3695, _d3696, _d3697, _d3698, _d3699}),
                    .FORW_LADDRAO({_d3700, _d3701, _d3702, _d3703, _d3704, _d3705, _d3706, _d3707, _d3708, _d3709, _d3710, _d3711, _d3712,
                   _d3713, _d3714, _d3715}),
                    .FORW_UADDRBO({_d3716, _d3717, _d3718, _d3719, _d3720, _d3721, _d3722, _d3723, _d3724, _d3725, _d3726, _d3727, _d3728,
                   _d3729, _d3730, _d3731}),
                    .FORW_LADDRBO({_d3732, _d3733, _d3734, _d3735, _d3736, _d3737, _d3738, _d3739, _d3740, _d3741, _d3742, _d3743, _d3744,
                   _d3745, _d3746, _d3747}),
                    .FORW_UA0CLKO(_d3748), .FORW_UA0ENO(_d3749), .FORW_UA0WEO(_d3750), .FORW_LA0CLKO(_d3751), .FORW_LA0ENO(_d3752),
                    .FORW_LA0WEO(_d3753), .FORW_UA1CLKO(_d3754), .FORW_UA1ENO(_d3755), .FORW_UA1WEO(_d3756), .FORW_LA1CLKO(_d3757),
                    .FORW_LA1ENO(_d3758), .FORW_LA1WEO(_d3759), .FORW_UB0CLKO(_d3760), .FORW_UB0ENO(_d3761), .FORW_UB0WEO(_d3762), .FORW_LB0CLKO(_d3763),
                    .FORW_LB0ENO(_d3764), .FORW_LB0WEO(_d3765), .FORW_UB1CLKO(_d3766), .FORW_UB1ENO(_d3767), .FORW_UB1WEO(_d3768), .FORW_LB1CLKO(_d3769),
                    .FORW_LB1ENO(_d3770), .FORW_LB1WEO(_d3771), .CLOCKA({_d3772, _d3773, _d3774, _d3775}),
                    .CLOCKB({_d3776, _d3777, _d3778, _d3779}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7452_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7454_10, na7455_9, na7456_10, na7458_9, na7459_10, na7460_9, na7462_10, na7463_9, na7464_10, na7466_9,
                   na7467_10, na7468_9, na7470_10, na7471_9, na7472_10, na7474_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7475_10, na7476_9, na7478_10, na7479_9, na7480_10,
                   na7482_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_01_80_00_00_00_00_03_03_00_00_00_23_03_13_23_00_00),
             .INIT_00(320'h22129e03b8e7fa9ef01cea789ff3c9003e0f24090271ce27890279c4f90761e07060f8a73c9e793c),
             .INIT_01(320'h0639c4a409f0129e27b8e7129ee39c4a4094a088003c04a789e6129025282213c001204fb9c4a528),
             .INIT_02(320'hf241c0701a0701a0700a43129411094f00000120e7fa8f7389ea5294a088003c04a789e831ce253d),
             .INIT_03(320'hea428ee389e753d4a05c47b9c4f79cea5294a504424004801c4ff9e48389ff3c90713fe7920e27fc),
             .INIT_04(320'he75214771c4f3a90a3b8e279d4851dc713cea428ee389e75214771c4f3a90a3b8e279d4851dc713c),
             .INIT_05(320'hef53dc73894813e0253c4f13ae73c9e5f9a4f7a9ee39c4a409e693cd27bd4a5294110948028ee389),
             .INIT_06(320'he693dea7b8e7129027c04a789e275ce7920fa054e693dea7b8e7129027c04a789e275ce793cbf349),
             .INIT_07(320'he03c94a50442520e039a4f7a9f0129e2789d739e4f3544a79a4f7a9027c04a789e275ce7920fa054),
             .INIT_08(320'h4f71ce253dc73894812941100e2928625044241da73dc06c09e753e41d8781c183a53ec5387e7d02),
             .INIT_09(320'h804284a5282238ad2549e27c04a7894714047b9ef7388f20094795ec25204a1104a5044001e0253c),
             .INIT_0A(320'he0b940e83c1683c10781e5021f603c08020e07c10f108e7b94c4f9a05213a48140c282002e015100),
             .INIT_0B(320'ha613c5753a4f149e279aa25384f12048108c22904a529411094a41c20000e7fb4f603c1711f0879f),
             .INIT_0C(320'h4f3c94a5282201cdf13e4f37c4f93cdf13e4f13f4a529411094f01cf8788fa53c5001b5291c5011e),
             .INIT_0D(320'h9d240a627cd028185040858360d101085094a5294a5294111c4a769e7b894ed3cf7129da79ee253f),
             .INIT_0E(320'h0f038a0681c682007b010f0200f03e0f03e08788473dca627cd021444d8a04281a52c10d108a5a90),
             .INIT_0F(320'h4a1284a504425294a5294a40027b81c0ba1e041c0f11f0879fe783cf07c1e7821e07140e02007b01),
             .INIT_10(320'h02b8000300e23e9c2bc9c2bc9c2bc9c2bc9c2bc9c2bc9c2bc9c2bc9423dcea79ff23dcea40847b9d),
             .INIT_11(320'h024085015c4abe9073fe47d3c0011e0253c4f39c4f11de75204810a0701c0681c0681c0681c0681c),
             .INIT_12(320'h4a504010044278afa400578094f13ca2758c27890241f4839ff23e9e0008f0129e279ce2788ef3a9),
             .INIT_13(320'h4f3800001cea79c073a9e739d4f39cea79ce753de713de0389ef01c4a52822120fa4c94a08807529),
             .INIT_14(320'he70004738047800f001e003c007800f001e003dc0753ee03a9f701d4f380e753cc701cea79c0039d),
             .INIT_15(320'h4f3c9f810802409f812941109e00090012002400480090713c027dc0752048398e491ce6288473a9),
             .INIT_16(320'h2213c0779c4a5282213c0001d41d8781c183831cf25004812002400480090013c401204f3c9e2b9e),
             .INIT_17(320'h3f3c0e039e0713f4069cf621c3f3c0a7b10e1f9e073d8a70fcf0389ff3c9e03f80793cf279e4a528),
             .INIT_18(320'h4a3bce25294a08848389ff3c9e275cc7a90e1f9e07920e27fcf2789d731ea4387e781e48389f629c),
             .INIT_19(320'he639e4f3a90279e4f50761e07060fe4a5282213cf23bce2529411090039fea51de71204d39ce7398),
             .INIT_1A(320'hf039fff95e073fff2bc0e7d40427e907b80ea79c073a9fa4004fd20f001f483c00739cea7e907800),
             .INIT_1B(320'h4a0884f000063804f120480094f50761e07060e9f8148e293b4e15f4781f483c0e7ffe5781cfffca),
             .INIT_1C(320'he73a9027880f11ce73a902788e739d4813c4739cea409e239ce75204f11ce73a902788fa79ce7529),
             .INIT_1D(320'h4f3dc4739cea409e7b88e739d4813cf711ce73a9027880f11de73a9027880f11ce73a9027880f11c),
             .INIT_1E(320'hd739e4f36ae693dea789d739e4f2fcd27bd4db9e5218941100e275ce793c57349ef5286250442400),
             .INIT_1F(320'he0389f8128ef3894a5044241f4992941100ea5294a08020088483e9e7b89fa79ee79294a50440389),
             .INIT_20(320'he03a9e701cea798e039d4f380073a9e70000039d4f380e753ce73a9e739d4f39cea7bce27bc0713d),
             .INIT_21(320'h023c007800f001e003c007800f001e003c007800f001e003c007800f001e003c007b80ea7dc0753e),
             .INIT_22(320'h3b0f038307f27a9c7368ef3890240048009001200241ee03a90241cc73e8e73144239d4ef800237c),
             .INIT_23(320'h4800900120024004f1004813cf27e0f25294a52941109e03a94779c4f790ef0fc3f0e0e1f89e27a8),
             .INIT_24(320'h442a9aa7bd482b54d21c671b0c0290aa6a9ef53fea7a9ea51de71200750761e07060e0c73c940120),
             .INIT_25(320'he73c9027e0f27a83b0f038307f27bd0013c4f13fe793b8c01cb839dea7a9ea6b54d21c671b0c0290),
             .INIT_26(320'h02780f2409e03b8a70fcf2409001294a0884f01de71294a0884a5294f0000750761e07060fe4f13a),
             .INIT_27(320'hea79ff639e4f7a9e7fdcd27bd48120e275ce79204f3dc4f3c902780f2409e2009e03c902780f2409),
             .INIT_28(320'h57d1e07b0957289d8d5fc715f4781ec2548c220c4a5282213c00120ea0ec3c0e0c1e90e7fd8e793d),
             .INIT_29(320'h4a1294a518441894a088483c007800f001e003c007800f00094a0880218941109483944ec6afe39c),
             .INIT_2A(320'hf001e003c007800f001e0011ee6d1ae7bdcc012047b9b46b98027e04a709c2529478094780947800),
             .INIT_2B(320'hf001e073a0f001e003c0e741e003c00781ce83200001cda798027c0001288252941109e2b4952789),
             .INIT_2C(320'h4279e4739c4a52822120073fd4a39ce2409a739ce73094739c4a5294110907800d2549e27c007800),
             .INIT_2D(320'h4813c40788e739d4813c4739cea409e239ce75204f11ce73a902788e739d4813c47d3ce73a94a504),
             .INIT_2E(320'he239ce75204f3dc4739cea409e7b88e739d4813c40788e739d4813c40788e739d4813c40788e739d),
             .INIT_2F(320'hf279b57349ef53c4eb9cf2797e693dea6dcf290c4a0880713ae73c9e2b9a4f7a943128221200279e),
             .INIT_30(320'h0251ce71294a52822120fa4c94a088075294a504010044241f4f3dc4fd3cf73c94a5282201c4eb9c),
             .INIT_31(320'he039d4ef1c073a9e7000e753ce0000073a9df01cea77ce753be73a9df39d4f39c4f380e279c0713f),
             .INIT_32(320'h024004800900120df00047780ea40906f1c9237cc5108e753be0008df008ef01d4f780ea7bc0753b),
             .INIT_33(320'h42780e73894a50442780ef0fc3f0e0e1c094a50442529e03bd48388e7389ef0fc3f0e0e1c0900120),
             .INIT_34(320'h4ff104728fe53bd4f7a9ef520e239ce2409e143dea41c4739c4f50761e07060e94a0094a5294a504),
             .INIT_35(320'hef53dea6b54d0140e2000701c0c31465228835a9ad53dea415aa690e03818628ca45106b535aa7bd),
             .INIT_36(320'he73984a39ce25294a0884a5294f01f0291c5710761e07060fec254047387e1f87070ec425294d6a9),
             .INIT_37(320'h02788df39d4813c46f9cea409e23e9df39d4a5282213cf239ce2529411090039fea51ce71204d39c),
             .INIT_38(320'he201c4739cea409e201c4739cea409e201c4739cea409e201c4739cea409e239ce75204f11ce73a9),
             .INIT_39(320'h6250440389d739e4f15cd27bd4a189411090013cf711be73a90279ee237ce75204f3dc46f9cea409),
             .INIT_3A(320'h4a52822120fa79ee27e9e7b9e4a52941100e275ce793cdab9a4f7a9e275ce793cbf349ef536e7948),
             .INIT_3B(320'he277c0713be71294a088483883b0f038307c514a52128f251e4ef98da789de39ff2789de39ff2789),
             .INIT_3C(320'he27984a788df389027e94ef80e277ce25294a50442789df3894fd3ce237ce253f4f388df3894a37c),
             .INIT_3D(320'h4a5294a13d424e94138de71adff09cc7b884111cc73c824310c410483310c320822120df389da529),
             .INIT_3E(320'hba5294a5294a529411094a53c480094a1082701b000004a786403e94a5294a000831094a50442409),
             .INIT_3F(320'h4a9294a5294a5294a528221284a5294a5294a474fa008180ec44180a308b8020ca100605f80a4188),
             .INIT_40(320'hc630cc0f7f66fe3f8fe31819cf0f9de73ff63e800000000000000003ff8ac212c6390c43800873e9),
             .INIT_41(320'h1f07f601808208000d8021ce4c02e0fe1e01006e6018c9b3e3e0d9fc0c1fe607ea10a367c78c621f),
             .INIT_42(320'h4a5205601e4b3f0f821038158027e847d8ce006c3b085fa1040179de5387b83ecff31f1fc63e0fe3),
             .INIT_43(320'h180401fd48fa91c1f0851fd442811f2010c00078b2f83181800b88529c9c1f064425094a5294a529),
             .INIT_44(320'h522f8bb000b0f83fa91f5f07c2147f010bf003ec42558027e06001807c001fd16e0f8b214a72707c),
             .INIT_45(320'hc310904090230866210c56009c7008f712956129027fc5801004044e2f8b07e84001985a917630c4),
             .INIT_46(320'h2701b000004a786403f44a500041884a528f8a0ac2009fab1e4f10cfab08027e84810b0700be2fea),
             .INIT_47(320'h001094a088481004a0884a5290015f4a504403804f0c807d280020c42529411094a529e241f4a10c),
             .INIT_48(320'hde390172e266f13d500810300e73602000803188431294a5044252048088031094a50442409f8000),
             .INIT_49(320'h40180bed63b100a462787f1e0641294a52907d8c4fc08400884a12aff9294310e5395f011094a409),
             .INIT_4A(320'h4a5e0b811f98060310e0f9838200020110021c0c032dbf079806c000297f79180060804009080180),
             .INIT_4B(320'h011295b9294a50071d2042928faf9cff2ffe9feb463f307800f9cde233e0fe10a87d60b91094a529),
             .INIT_4C(320'h0011044100473f68600806380feb94f8e9cff4fc1d3eb04fe4425294a529027e0983fc07d9f5bd8b),
             .INIT_4D(320'h4a48053d2042928fad14fef9ac7d08f8c1a785f4b638f04002fa1fc533e0f8240e4b886308002c1b),
             .INIT_4E(320'he7f50401004701fd7c7cff21cff4fc1c3eb05fe4425294a529027e0b83fc07e9f3dd87031295b929),
             .INIT_4F(320'h411ec00008021ea60000024090500f5300000200040147a9800001002c10a020c241873820482004),
             .INIT_50(320'h48383511002230a03a904a5294a49c621295cd2902128f9c857a19280be80209077c1f183c063100),
             .INIT_51(320'h4812047c106b7f0c5198a41094a5294a528221244a5294a52948109022082019e250060607c40920),
             .INIT_52(320'hfc2805a84802000c7dad67c0402100a7d40a35bf663f4fa28d6fd14c2014833e0cb704425094a529),
             .INIT_53(320'h80b184dd17102a08fe90bf0405ed18f2810ba8081029f060004100840290fabe2470008400d6fd98),
             .INIT_54(320'h423094804002340e00000014042529423ed6fc0800300063e020108053eafa0404701f5ec1c13314),
             .INIT_55(320'h02808203ffe03fcd8008f005c0110846009488004681c001094a10407ffc07f9b0011e00b802212b),
             .INIT_56(320'h470144a088c115c07960fb01f0025c0601bb0140413e8e110902b80d2c09da0002218006c12073f6),
             .INIT_57(320'h423e02230b023e09fbdec67f8f633fc7b19faa95b2088c02089fbc8c033fa7a00a57f8f4018cff0a),
             .INIT_58(320'he579964280380fd07407fd4806b538ff1bc88008040073f404c6f9ba54fff3118f9380411094a7e9),
             .INIT_59(320'hc920dc6300c6707a64130c33004c3fa34040a33d0009804495d7f98c0311c02bb007f9ff32df4324),
             .INIT_5A(320'hdf79c4006122009fa5083a3e0262a0e809cf84884f3e10240c41f9c3f407ef4fd0741d0741fe9c90),
             .INIT_5B(320'hfbdc83843f4a5083fff0e7fcc0fc60e73a44291f011094a5294808700060085294a52947c041907c),
             .INIT_5C(320'h0000004010043ec3fd083a53f73107e879fce03d0839fce03d08321f7018d83a1e803f400ec3f3e1),
             .INIT_5D(320'h318c6318c6318c6002d6b5ad6b5ad6b5ad6000c6318c6318c6318c6000c6318c6318c6318c600000),
             .INIT_5E(320'h739ce739ce739ce000c6318c6318c6318c6002d6b5ad6b5ad6b5ad6001ce739ce739ce739ce000c6),
             .INIT_5F(320'h0000042108421084000000000421084210840000000004421084210002d6b5ad6b5ad6b5ad6001ce),
             .INIT_60(320'hd8c711ce6b1ee2358c635ee605ae6b58240cae6302c0242108421084210842108400000000040000),
             .INIT_61(320'h1847318b7b580731847318f6b08c2b0ec7b1ed619846a580225813352c09d8f295a6239cd631ac63),
             .INIT_62(320'h5815b1c5631ed63dac121cc3b98c0bd817b5ec6b00000000000000000000000230ac3b1ab7b58073),
             .INIT_63(320'h089421401f18c6008c735cd63182409ef43181735ec120652b98c0b0044a1080a048631aa6318d53),
             .INIT_64(320'h821100a06b5857304e600000000000900615cc60580225084010442104411692a088121e57318160),
             .INIT_65(320'h9af23dac72de47b5ad231cf6b0687198e6302f6318a6b042139cf39048735cc7a18d7b5ad6302529),
             .INIT_66(320'h1ac4b18d3b1ac63581720a52352f2b08d6bd823b8a56b1ad791ad7b02f2302d2300161d8e6b1cd4b),
             .INIT_67(320'h88262eb3eeca36a35c9514c1177d9d56d19b9aa498a20fbbacdab28048635cc6358c121cd6358e63),
             .INIT_68(320'ha92e6ca36aeb3ee14c1135c9556d1977d9d98a20b9aa4dab28fbbac254d704453675df4655ba92e6),
             .INIT_69(320'h290842002000c63194a4210805ce2b5a56090e635ae6302d4302d6304453254d74655b675df88262),
             .INIT_6A(320'h1ce631ac72420000487358d6b5cc605c66bdc56b1ab60802008002000c63194a4210800800318c65),
             .INIT_6B(320'h94a5bda94092a5bda84012a5bdab40d4952ded52925719ed6a00d7bca54200c73da81318c5a9816b),
             .INIT_6C(320'h01063000631ad639882ad0c4a02d631c94012a6b4a86b9ad718c5731ac4a50803da67a5027b1892a),
             .INIT_6D(320'h31800318c6318c6318c6318842000008c1bd803bdec120656b1ce731cc015856bdc46b1800000000),
             .INIT_6E(320'hb5800739ce739ce739ce73800318c6318c6318c631800b5ad6b5ad6b5ad6b5800318c6318c6318c6),
             .INIT_6F(320'h84000b5ad6b5ad6b5ad6b5800739ce739ce739ce73800318c6318c6318c631800b5ad6b5ad6b5ad6),
             .INIT_70(320'h42108421084210000000001000000000108421084210000000001084210842100000000011084210),
             .INIT_71(320'h00c3b948715ee615ef7302e6b9ee61d8d619802b0ad7b88d6398c730486358b73181600ad0842108),
             .INIT_72(320'h2940006c4b00c291c4415cd211c54952c1bd80295cc0ad8e609032b58e3b98c0b98c73294800037b),
             .INIT_73(320'h318c6318c6000219ac63de9430244158f2a18123509430466a1807300c1118d791ae335ce6300565),
             .INIT_74(320'h00000000000000000000000000000000000018d800000318c6318c6318c6318c6318c6318c6318c6),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6643 ( .DOA({_d3780, _d3781, _d3782, _d3783, _d3784, _d3785, _d3786, _d3787, _d3788, _d3789, _d3790, _d3791, _d3792, _d3793,
                   _d3794, _d3795, _d3796, _d3797, _d3798, _d3799, _d3800, _d3801, _d3802, _d3803, _d3804, _d3805, _d3806, _d3807, _d3808,
                   _d3809, _d3810, _d3811, _d3812, _d3813, _d3814, na6643_36, na6643_37, na6643_38, na6643_39, na6643_40}),
                    .DOAX({_d3815, _d3816, _d3817, _d3818, _d3819, _d3820, _d3821, _d3822, _d3823, _d3824, _d3825, _d3826, _d3827, _d3828,
                   _d3829, _d3830, _d3831, _d3832, _d3833, _d3834, _d3835, _d3836, _d3837, _d3838, _d3839, _d3840, _d3841, _d3842, _d3843,
                   _d3844, _d3845, _d3846, _d3847, _d3848, _d3849, _d3850, _d3851, _d3852, _d3853, _d3854}),
                    .DOB({_d3855, _d3856, _d3857, _d3858, _d3859, _d3860, _d3861, _d3862, _d3863, _d3864, _d3865, _d3866, _d3867, _d3868,
                   _d3869, _d3870, _d3871, _d3872, _d3873, _d3874, _d3875, _d3876, _d3877, _d3878, _d3879, _d3880, _d3881, _d3882, _d3883,
                   _d3884, _d3885, _d3886, _d3887, _d3888, _d3889, _d3890, _d3891, _d3892, _d3893, _d3894}),
                    .DOBX({_d3895, _d3896, _d3897, _d3898, _d3899, _d3900, _d3901, _d3902, _d3903, _d3904, _d3905, _d3906, _d3907, _d3908,
                   _d3909, _d3910, _d3911, _d3912, _d3913, _d3914, _d3915, _d3916, _d3917, _d3918, _d3919, _d3920, _d3921, _d3922, _d3923,
                   _d3924, _d3925, _d3926, _d3927, _d3928, _d3929, _d3930, _d3931, _d3932, _d3933, _d3934}),
                    .ECC1B_ERRA({_d3935, _d3936, _d3937, _d3938}),
                    .ECC1B_ERRB({_d3939, _d3940, _d3941, _d3942}),
                    .ECC2B_ERRA({_d3943, _d3944, _d3945, _d3946}),
                    .ECC2B_ERRB({_d3947, _d3948, _d3949, _d3950}),
                    .FORW_CAS_WRAO(_d3951), .FORW_CAS_WRBO(_d3952), .FORW_CAS_BMAO(_d3953), .FORW_CAS_BMBO(_d3954), .FORW_CAS_RDAO(_d3955),
                    .FORW_CAS_RDBO(_d3956), .FORW_UADDRAO({_d3957, _d3958, _d3959, _d3960, _d3961, _d3962, _d3963, _d3964, _d3965, _d3966,
                   _d3967, _d3968, _d3969, _d3970, _d3971, _d3972}),
                    .FORW_LADDRAO({_d3973, _d3974, _d3975, _d3976, _d3977, _d3978, _d3979, _d3980, _d3981, _d3982, _d3983, _d3984, _d3985,
                   _d3986, _d3987, _d3988}),
                    .FORW_UADDRBO({_d3989, _d3990, _d3991, _d3992, _d3993, _d3994, _d3995, _d3996, _d3997, _d3998, _d3999, _d4000, _d4001,
                   _d4002, _d4003, _d4004}),
                    .FORW_LADDRBO({_d4005, _d4006, _d4007, _d4008, _d4009, _d4010, _d4011, _d4012, _d4013, _d4014, _d4015, _d4016, _d4017,
                   _d4018, _d4019, _d4020}),
                    .FORW_UA0CLKO(_d4021), .FORW_UA0ENO(_d4022), .FORW_UA0WEO(_d4023), .FORW_LA0CLKO(_d4024), .FORW_LA0ENO(_d4025),
                    .FORW_LA0WEO(_d4026), .FORW_UA1CLKO(_d4027), .FORW_UA1ENO(_d4028), .FORW_UA1WEO(_d4029), .FORW_LA1CLKO(_d4030),
                    .FORW_LA1ENO(_d4031), .FORW_LA1WEO(_d4032), .FORW_UB0CLKO(_d4033), .FORW_UB0ENO(_d4034), .FORW_UB0WEO(_d4035), .FORW_LB0CLKO(_d4036),
                    .FORW_LB0ENO(_d4037), .FORW_LB0WEO(_d4038), .FORW_UB1CLKO(_d4039), .FORW_UB1ENO(_d4040), .FORW_UB1WEO(_d4041), .FORW_LB1CLKO(_d4042),
                    .FORW_LB1ENO(_d4043), .FORW_LB1WEO(_d4044), .CLOCKA({_d4045, _d4046, _d4047, _d4048}),
                    .CLOCKB({_d4049, _d4050, _d4051, _d4052}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7498_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7499_10, na7500_9, na7502_10, na7503_9, na7504_10, na7506_9, na7507_10, na7508_9, na7510_10, na7511_9,
                   na7512_10, na7514_9, na7515_10, na7516_9, na7518_10, na7519_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7520_10, na7522_9, na7523_10, na7524_9, na7526_10,
                   na7527_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_02_80_15_00_00_00_03_03_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6644 ( .DOA({_d4053, _d4054, _d4055, _d4056, _d4057, _d4058, _d4059, _d4060, _d4061, _d4062, _d4063, _d4064, _d4065, _d4066,
                   _d4067, _d4068, _d4069, _d4070, _d4071, _d4072, na6644_21, na6644_22, na6644_23, na6644_24, na6644_25, na6644_26,
                   na6644_27, na6644_28, na6644_29, na6644_30, na6644_31, na6644_32, na6644_33, na6644_34, na6644_35, na6644_36, na6644_37,
                   na6644_38, na6644_39, na6644_40}),
                    .DOAX({_d4073, _d4074, _d4075, _d4076, _d4077, _d4078, _d4079, _d4080, _d4081, _d4082, _d4083, _d4084, _d4085, _d4086,
                   _d4087, _d4088, _d4089, _d4090, _d4091, _d4092, _d4093, _d4094, _d4095, _d4096, _d4097, _d4098, _d4099, _d4100, _d4101,
                   _d4102, _d4103, _d4104, _d4105, _d4106, _d4107, _d4108, _d4109, _d4110, _d4111, _d4112}),
                    .DOB({_d4113, _d4114, _d4115, _d4116, _d4117, _d4118, _d4119, _d4120, _d4121, _d4122, _d4123, _d4124, _d4125, _d4126,
                   _d4127, _d4128, _d4129, _d4130, _d4131, _d4132, _d4133, _d4134, _d4135, _d4136, _d4137, _d4138, _d4139, _d4140, _d4141,
                   _d4142, _d4143, _d4144, _d4145, _d4146, _d4147, _d4148, _d4149, _d4150, _d4151, _d4152}),
                    .DOBX({_d4153, _d4154, _d4155, _d4156, _d4157, _d4158, _d4159, _d4160, _d4161, _d4162, _d4163, _d4164, _d4165, _d4166,
                   _d4167, _d4168, _d4169, _d4170, _d4171, _d4172, _d4173, _d4174, _d4175, _d4176, _d4177, _d4178, _d4179, _d4180, _d4181,
                   _d4182, _d4183, _d4184, _d4185, _d4186, _d4187, _d4188, _d4189, _d4190, _d4191, _d4192}),
                    .ECC1B_ERRA({_d4193, _d4194, _d4195, _d4196}),
                    .ECC1B_ERRB({_d4197, _d4198, _d4199, _d4200}),
                    .ECC2B_ERRA({_d4201, _d4202, _d4203, _d4204}),
                    .ECC2B_ERRB({_d4205, _d4206, _d4207, _d4208}),
                    .FORW_CAS_WRAO(_d4209), .FORW_CAS_WRBO(_d4210), .FORW_CAS_BMAO(_d4211), .FORW_CAS_BMBO(_d4212), .FORW_CAS_RDAO(_d4213),
                    .FORW_CAS_RDBO(_d4214), .FORW_UADDRAO({_d4215, _d4216, _d4217, _d4218, _d4219, _d4220, _d4221, _d4222, _d4223, _d4224,
                   _d4225, _d4226, _d4227, _d4228, _d4229, _d4230}),
                    .FORW_LADDRAO({_d4231, _d4232, _d4233, _d4234, _d4235, _d4236, _d4237, _d4238, _d4239, _d4240, _d4241, _d4242, _d4243,
                   _d4244, _d4245, _d4246}),
                    .FORW_UADDRBO({_d4247, _d4248, _d4249, _d4250, _d4251, _d4252, _d4253, _d4254, _d4255, _d4256, _d4257, _d4258, _d4259,
                   _d4260, _d4261, _d4262}),
                    .FORW_LADDRBO({_d4263, _d4264, _d4265, _d4266, _d4267, _d4268, _d4269, _d4270, _d4271, _d4272, _d4273, _d4274, _d4275,
                   _d4276, _d4277, _d4278}),
                    .FORW_UA0CLKO(_d4279), .FORW_UA0ENO(_d4280), .FORW_UA0WEO(_d4281), .FORW_LA0CLKO(_d4282), .FORW_LA0ENO(_d4283),
                    .FORW_LA0WEO(_d4284), .FORW_UA1CLKO(_d4285), .FORW_UA1ENO(_d4286), .FORW_UA1WEO(_d4287), .FORW_LA1CLKO(_d4288),
                    .FORW_LA1ENO(_d4289), .FORW_LA1WEO(_d4290), .FORW_UB0CLKO(_d4291), .FORW_UB0ENO(_d4292), .FORW_UB0WEO(_d4293), .FORW_LB0CLKO(_d4294),
                    .FORW_LB0ENO(_d4295), .FORW_LB0WEO(_d4296), .FORW_UB1CLKO(_d4297), .FORW_UB1ENO(_d4298), .FORW_UB1WEO(_d4299), .FORW_LB1CLKO(_d4300),
                    .FORW_LB1ENO(_d4301), .FORW_LB1WEO(_d4302), .CLOCKA({_d4303, _d4304, _d4305, _d4306}),
                    .CLOCKB({_d4307, _d4308, _d4309, _d4310}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7535_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, na7536_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7538_10, na7539_9, na7540_10, na7542_9, na7543_10, na7544_9, na7546_10, na7547_9, na7548_10, na7550_9,
                   na7551_10, na7552_9, na7554_10, na7555_9, na7556_10, na7558_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7559_9, 1'b1, na7560_9, na7562_10, na7563_9, na7564_10,
                   na7566_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na7567_10, na7568_9, na7570_10, na7571_9, na7572_10, na7574_9, na7575_10, na7576_9, na7578_10, na7579_9,
                   na7580_10, na7582_9, na7583_10, na7584_9, na7586_10, na7587_9, na7588_10, na7590_9, na7591_10, na7592_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na7602_10, na7603_9, na7604_10, na7606_9, na7607_10, na7608_9, na7618_10, na7619_9, na7620_10, na7624_9,
                   na7625_10, na7626_9, na7631_10, na7634_9, na7635_10, na7636_9, na7638_10, na7639_9, na7640_10, na7642_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_00_16_80_B5_03_03_00_03_03_00_00_13_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6645 ( .DOA({na6645_1, na6645_2, na6645_3, na6645_4, na6645_5, na6645_6, na6645_7, na6645_8, na6645_9, na6645_10, na6645_11,
                   na6645_12, na6645_13, na6645_14, na6645_15, na6645_16, na6645_17, na6645_18, na6645_19, na6645_20, na6645_21, na6645_22,
                   na6645_23, na6645_24, na6645_25, na6645_26, na6645_27, na6645_28, na6645_29, na6645_30, na6645_31, na6645_32, na6645_33,
                   na6645_34, na6645_35, na6645_36, na6645_37, na6645_38, na6645_39, na6645_40}),
                    .DOAX({_d4311, _d4312, _d4313, _d4314, _d4315, _d4316, _d4317, _d4318, _d4319, _d4320, _d4321, _d4322, _d4323, _d4324,
                   _d4325, _d4326, _d4327, _d4328, _d4329, _d4330, _d4331, _d4332, _d4333, _d4334, _d4335, _d4336, _d4337, _d4338, _d4339,
                   _d4340, _d4341, _d4342, _d4343, _d4344, _d4345, _d4346, _d4347, _d4348, _d4349, _d4350}),
                    .DOB({_d4351, _d4352, _d4353, _d4354, _d4355, _d4356, _d4357, _d4358, _d4359, _d4360, _d4361, _d4362, _d4363, _d4364,
                   _d4365, _d4366, _d4367, _d4368, _d4369, _d4370, _d4371, _d4372, _d4373, _d4374, _d4375, _d4376, _d4377, _d4378, _d4379,
                   _d4380, _d4381, _d4382, _d4383, _d4384, _d4385, _d4386, _d4387, _d4388, _d4389, _d4390}),
                    .DOBX({_d4391, _d4392, _d4393, _d4394, _d4395, _d4396, _d4397, _d4398, _d4399, _d4400, _d4401, _d4402, _d4403, _d4404,
                   _d4405, _d4406, _d4407, _d4408, _d4409, _d4410, _d4411, _d4412, _d4413, _d4414, _d4415, _d4416, _d4417, _d4418, _d4419,
                   _d4420, _d4421, _d4422, _d4423, _d4424, _d4425, _d4426, _d4427, _d4428, _d4429, _d4430}),
                    .ECC1B_ERRA({_d4431, _d4432, _d4433, _d4434}),
                    .ECC1B_ERRB({_d4435, _d4436, _d4437, _d4438}),
                    .ECC2B_ERRA({_d4439, _d4440, _d4441, _d4442}),
                    .ECC2B_ERRB({_d4443, _d4444, _d4445, _d4446}),
                    .FORW_CAS_WRAO(_d4447), .FORW_CAS_WRBO(_d4448), .FORW_CAS_BMAO(_d4449), .FORW_CAS_BMBO(_d4450), .FORW_CAS_RDAO(_d4451),
                    .FORW_CAS_RDBO(_d4452), .FORW_UADDRAO({_d4453, _d4454, _d4455, _d4456, _d4457, _d4458, _d4459, _d4460, _d4461, _d4462,
                   _d4463, _d4464, _d4465, _d4466, _d4467, _d4468}),
                    .FORW_LADDRAO({_d4469, _d4470, _d4471, _d4472, _d4473, _d4474, _d4475, _d4476, _d4477, _d4478, _d4479, _d4480, _d4481,
                   _d4482, _d4483, _d4484}),
                    .FORW_UADDRBO({_d4485, _d4486, _d4487, _d4488, _d4489, _d4490, _d4491, _d4492, _d4493, _d4494, _d4495, _d4496, _d4497,
                   _d4498, _d4499, _d4500}),
                    .FORW_LADDRBO({_d4501, _d4502, _d4503, _d4504, _d4505, _d4506, _d4507, _d4508, _d4509, _d4510, _d4511, _d4512, _d4513,
                   _d4514, _d4515, _d4516}),
                    .FORW_UA0CLKO(_d4517), .FORW_UA0ENO(_d4518), .FORW_UA0WEO(_d4519), .FORW_LA0CLKO(_d4520), .FORW_LA0ENO(_d4521),
                    .FORW_LA0WEO(_d4522), .FORW_UA1CLKO(_d4523), .FORW_UA1ENO(_d4524), .FORW_UA1WEO(_d4525), .FORW_LA1CLKO(_d4526),
                    .FORW_LA1ENO(_d4527), .FORW_LA1WEO(_d4528), .FORW_UB0CLKO(_d4529), .FORW_UB0ENO(_d4530), .FORW_UB0WEO(_d4531), .FORW_LB0CLKO(_d4532),
                    .FORW_LB0ENO(_d4533), .FORW_LB0WEO(_d4534), .FORW_UB1CLKO(_d4535), .FORW_UB1ENO(_d4536), .FORW_UB1WEO(_d4537), .FORW_LB1CLKO(_d4538),
                    .FORW_LB1ENO(_d4539), .FORW_LB1WEO(_d4540), .CLOCKA({_d4541, _d4542, _d4543, _d4544}),
                    .CLOCKB({_d4545, _d4546, _d4547, _d4548}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, na7643_9, 1'b1, na7644_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na7646_10, 1'b1, na7647_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7648_10, na7650_9, na7651_10, na7652_9, na7654_10, na7655_9, na7656_10, na7658_9, na7659_10, na7660_9,
                   na7710_10, na7711_9, na7712_10, na7714_9, na7715_10, na7716_9}),
                    .ADDRA1({na7717_10, na7718_9, na7719_10, na7720_9, na7721_10, na7722_9, na7724_10, na7725_9, na7726_10, na7731_9,
                   na7734_10, na7739_9, na7742_10, na7744_9, na7750_10, na7752_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7758_9, 1'b1, na7760_9, na7766_10, na7768_9, na7777_10,
                   na7779_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na7783_9, 1'b1, na7785_9, na7789_10, na7791_9, na7795_10,
                   na7797_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na7801_10, na7803_9, na7807_10, na7809_9, na7813_10, na7815_9, na7819_10, na7821_9, na7827_10, na7831_9, na7835_10,
                   na7839_9, na7843_10, na7847_9, na7851_10, na7855_9, na7859_10, na7863_9, na7867_10, na7871_9, na7875_10, na7879_9,
                   na7883_10, na7887_9, na7892_10, na7894_9, na7896_10, na7898_9, na7900_10, na7902_9, na7904_10, na7906_9, na7907_10,
                   na7908_9, na7909_10, na7911_9, na7913_10, na7914_9, na7915_10, na7916_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na7917_10, na7919_9, na7920_10, na7921_9, na7923_10, na7925_9, na7927_10, na7929_9, na7931_10, na7932_9, na7933_10,
                   na7935_9, na7937_10, na7939_9, na7941_10, na7943_9, na7945_10, na7946_9, na7947_10, na7949_9, na7951_10, na7956_9,
                   na7958_10, na7960_9, na7962_10, na7964_9, na7965_10, na7968_9, na7969_10, na7970_9, na7972_10, na7973_9, na7974_10,
                   na7976_9, na7977_10, na7978_9, na7980_10, na7981_9, na7982_10, na7984_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_///AND/      x59y65     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6646_4 ( .OUT(na6646_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2519_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6646_6 ( .RAM_O2(na6646_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6646_2), .COMP_OUT(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_02_80_15_00_00_00_03_03_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6647 ( .DOA({_d4549, _d4550, _d4551, _d4552, _d4553, _d4554, _d4555, _d4556, _d4557, _d4558, _d4559, _d4560, _d4561, _d4562,
                   _d4563, _d4564, _d4565, _d4566, _d4567, _d4568, na6647_21, na6647_22, na6647_23, na6647_24, na6647_25, na6647_26,
                   na6647_27, na6647_28, na6647_29, na6647_30, na6647_31, na6647_32, na6647_33, na6647_34, na6647_35, na6647_36, na6647_37,
                   na6647_38, na6647_39, na6647_40}),
                    .DOAX({_d4569, _d4570, _d4571, _d4572, _d4573, _d4574, _d4575, _d4576, _d4577, _d4578, _d4579, _d4580, _d4581, _d4582,
                   _d4583, _d4584, _d4585, _d4586, _d4587, _d4588, _d4589, _d4590, _d4591, _d4592, _d4593, _d4594, _d4595, _d4596, _d4597,
                   _d4598, _d4599, _d4600, _d4601, _d4602, _d4603, _d4604, _d4605, _d4606, _d4607, _d4608}),
                    .DOB({_d4609, _d4610, _d4611, _d4612, _d4613, _d4614, _d4615, _d4616, _d4617, _d4618, _d4619, _d4620, _d4621, _d4622,
                   _d4623, _d4624, _d4625, _d4626, _d4627, _d4628, _d4629, _d4630, _d4631, _d4632, _d4633, _d4634, _d4635, _d4636, _d4637,
                   _d4638, _d4639, _d4640, _d4641, _d4642, _d4643, _d4644, _d4645, _d4646, _d4647, _d4648}),
                    .DOBX({_d4649, _d4650, _d4651, _d4652, _d4653, _d4654, _d4655, _d4656, _d4657, _d4658, _d4659, _d4660, _d4661, _d4662,
                   _d4663, _d4664, _d4665, _d4666, _d4667, _d4668, _d4669, _d4670, _d4671, _d4672, _d4673, _d4674, _d4675, _d4676, _d4677,
                   _d4678, _d4679, _d4680, _d4681, _d4682, _d4683, _d4684, _d4685, _d4686, _d4687, _d4688}),
                    .ECC1B_ERRA({_d4689, _d4690, _d4691, _d4692}),
                    .ECC1B_ERRB({_d4693, _d4694, _d4695, _d4696}),
                    .ECC2B_ERRA({_d4697, _d4698, _d4699, _d4700}),
                    .ECC2B_ERRB({_d4701, _d4702, _d4703, _d4704}),
                    .FORW_CAS_WRAO(_d4705), .FORW_CAS_WRBO(_d4706), .FORW_CAS_BMAO(_d4707), .FORW_CAS_BMBO(_d4708), .FORW_CAS_RDAO(_d4709),
                    .FORW_CAS_RDBO(_d4710), .FORW_UADDRAO({_d4711, _d4712, _d4713, _d4714, _d4715, _d4716, _d4717, _d4718, _d4719, _d4720,
                   _d4721, _d4722, _d4723, _d4724, _d4725, _d4726}),
                    .FORW_LADDRAO({_d4727, _d4728, _d4729, _d4730, _d4731, _d4732, _d4733, _d4734, _d4735, _d4736, _d4737, _d4738, _d4739,
                   _d4740, _d4741, _d4742}),
                    .FORW_UADDRBO({_d4743, _d4744, _d4745, _d4746, _d4747, _d4748, _d4749, _d4750, _d4751, _d4752, _d4753, _d4754, _d4755,
                   _d4756, _d4757, _d4758}),
                    .FORW_LADDRBO({_d4759, _d4760, _d4761, _d4762, _d4763, _d4764, _d4765, _d4766, _d4767, _d4768, _d4769, _d4770, _d4771,
                   _d4772, _d4773, _d4774}),
                    .FORW_UA0CLKO(_d4775), .FORW_UA0ENO(_d4776), .FORW_UA0WEO(_d4777), .FORW_LA0CLKO(_d4778), .FORW_LA0ENO(_d4779),
                    .FORW_LA0WEO(_d4780), .FORW_UA1CLKO(_d4781), .FORW_UA1ENO(_d4782), .FORW_UA1WEO(_d4783), .FORW_LA1CLKO(_d4784),
                    .FORW_LA1ENO(_d4785), .FORW_LA1WEO(_d4786), .FORW_UB0CLKO(_d4787), .FORW_UB0ENO(_d4788), .FORW_UB0WEO(_d4789), .FORW_LB0CLKO(_d4790),
                    .FORW_LB0ENO(_d4791), .FORW_LB0WEO(_d4792), .FORW_UB1CLKO(_d4793), .FORW_UB1ENO(_d4794), .FORW_UB1WEO(_d4795), .FORW_LB1CLKO(_d4796),
                    .FORW_LB1ENO(_d4797), .FORW_LB1WEO(_d4798), .CLOCKA({_d4799, _d4800, _d4801, _d4802}),
                    .CLOCKB({_d4803, _d4804, _d4805, _d4806}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na7985_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, na7986_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na7988_10, na7989_9, na7990_10, na7991_9, na7992_10, na7993_9, na7995_10, na7996_9, na7998_10, na7999_9,
                   na8001_10, na8002_9, na8004_10, na8005_9, na8007_10, na8008_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8010_9, 1'b1, na8011_9, na8013_10, na8014_9, na8016_10,
                   na8017_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na8019_10, na8020_9, na8022_10, na8023_9, na8025_10, na8026_9, na8028_10, na8029_9, na8031_10, na8032_9,
                   na8034_10, na8035_9, na8037_10, na8038_9, na8040_10, na8041_9, na8042_10, na8043_9, na8044_10, na8045_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na8046_10, na8047_9, na8048_10, na8049_9, na8050_10, na8051_9, na8052_10, na8053_9, na8054_10, na8055_9,
                   na8056_10, na8057_9, na8059_10, na8060_9, na8062_10, na8064_9, na8066_10, na8068_9, na8071_10, na8074_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_00_16_80_B5_03_03_00_03_03_00_00_13_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6648 ( .DOA({na6648_1, na6648_2, na6648_3, na6648_4, na6648_5, na6648_6, na6648_7, na6648_8, na6648_9, na6648_10, na6648_11,
                   na6648_12, na6648_13, na6648_14, na6648_15, na6648_16, na6648_17, na6648_18, na6648_19, na6648_20, na6648_21, na6648_22,
                   na6648_23, na6648_24, na6648_25, na6648_26, na6648_27, na6648_28, na6648_29, na6648_30, na6648_31, na6648_32, na6648_33,
                   na6648_34, na6648_35, na6648_36, na6648_37, na6648_38, na6648_39, na6648_40}),
                    .DOAX({_d4807, _d4808, _d4809, _d4810, _d4811, _d4812, _d4813, _d4814, _d4815, _d4816, _d4817, _d4818, _d4819, _d4820,
                   _d4821, _d4822, _d4823, _d4824, _d4825, _d4826, _d4827, _d4828, _d4829, _d4830, _d4831, _d4832, _d4833, _d4834, _d4835,
                   _d4836, _d4837, _d4838, _d4839, _d4840, _d4841, _d4842, _d4843, _d4844, _d4845, _d4846}),
                    .DOB({_d4847, _d4848, _d4849, _d4850, _d4851, _d4852, _d4853, _d4854, _d4855, _d4856, _d4857, _d4858, _d4859, _d4860,
                   _d4861, _d4862, _d4863, _d4864, _d4865, _d4866, _d4867, _d4868, _d4869, _d4870, _d4871, _d4872, _d4873, _d4874, _d4875,
                   _d4876, _d4877, _d4878, _d4879, _d4880, _d4881, _d4882, _d4883, _d4884, _d4885, _d4886}),
                    .DOBX({_d4887, _d4888, _d4889, _d4890, _d4891, _d4892, _d4893, _d4894, _d4895, _d4896, _d4897, _d4898, _d4899, _d4900,
                   _d4901, _d4902, _d4903, _d4904, _d4905, _d4906, _d4907, _d4908, _d4909, _d4910, _d4911, _d4912, _d4913, _d4914, _d4915,
                   _d4916, _d4917, _d4918, _d4919, _d4920, _d4921, _d4922, _d4923, _d4924, _d4925, _d4926}),
                    .ECC1B_ERRA({_d4927, _d4928, _d4929, _d4930}),
                    .ECC1B_ERRB({_d4931, _d4932, _d4933, _d4934}),
                    .ECC2B_ERRA({_d4935, _d4936, _d4937, _d4938}),
                    .ECC2B_ERRB({_d4939, _d4940, _d4941, _d4942}),
                    .FORW_CAS_WRAO(_d4943), .FORW_CAS_WRBO(_d4944), .FORW_CAS_BMAO(_d4945), .FORW_CAS_BMBO(_d4946), .FORW_CAS_RDAO(_d4947),
                    .FORW_CAS_RDBO(_d4948), .FORW_UADDRAO({_d4949, _d4950, _d4951, _d4952, _d4953, _d4954, _d4955, _d4956, _d4957, _d4958,
                   _d4959, _d4960, _d4961, _d4962, _d4963, _d4964}),
                    .FORW_LADDRAO({_d4965, _d4966, _d4967, _d4968, _d4969, _d4970, _d4971, _d4972, _d4973, _d4974, _d4975, _d4976, _d4977,
                   _d4978, _d4979, _d4980}),
                    .FORW_UADDRBO({_d4981, _d4982, _d4983, _d4984, _d4985, _d4986, _d4987, _d4988, _d4989, _d4990, _d4991, _d4992, _d4993,
                   _d4994, _d4995, _d4996}),
                    .FORW_LADDRBO({_d4997, _d4998, _d4999, _d5000, _d5001, _d5002, _d5003, _d5004, _d5005, _d5006, _d5007, _d5008, _d5009,
                   _d5010, _d5011, _d5012}),
                    .FORW_UA0CLKO(_d5013), .FORW_UA0ENO(_d5014), .FORW_UA0WEO(_d5015), .FORW_LA0CLKO(_d5016), .FORW_LA0ENO(_d5017),
                    .FORW_LA0WEO(_d5018), .FORW_UA1CLKO(_d5019), .FORW_UA1ENO(_d5020), .FORW_UA1WEO(_d5021), .FORW_LA1CLKO(_d5022),
                    .FORW_LA1ENO(_d5023), .FORW_LA1WEO(_d5024), .FORW_UB0CLKO(_d5025), .FORW_UB0ENO(_d5026), .FORW_UB0WEO(_d5027), .FORW_LB0CLKO(_d5028),
                    .FORW_LB0ENO(_d5029), .FORW_LB0WEO(_d5030), .FORW_UB1CLKO(_d5031), .FORW_UB1ENO(_d5032), .FORW_UB1WEO(_d5033), .FORW_LB1CLKO(_d5034),
                    .FORW_LB1ENO(_d5035), .FORW_LB1WEO(_d5036), .CLOCKA({_d5037, _d5038, _d5039, _d5040}),
                    .CLOCKB({_d5041, _d5042, _d5043, _d5044}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, na8079_9, 1'b1, na8082_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na8083_10, 1'b1, na8084_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na8086_10, na8088_9, na8090_10, na8100_9, na8102_10, na8105_9, na8108_10, na8110_9, na8112_10, na8114_9,
                   na8115_10, na8117_9, na8120_10, na8122_9, na8124_10, na8126_9}),
                    .ADDRA1({na8127_10, na8128_9, na8129_10, na8131_9, na8133_10, na8135_9, na8136_10, na8138_9, na8139_10, na8140_9,
                   na8141_10, na8143_9, na8144_10, na8145_9, na8146_10, na8147_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8148_9, 1'b1, na8149_9, na8150_10, na8153_9, na8155_10,
                   na8156_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8157_9, 1'b1, na8159_9, na8160_10, na8161_9, na8162_10,
                   na8163_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na8164_10, na8165_9, na8168_10, na8169_9, na8170_10, na8171_9, na8172_10, na8178_9, na8179_10, na8180_9, na8181_10,
                   na8188_9, na8189_10, na8191_9, na8193_10, na8194_9, na8195_10, na8196_9, na8198_10, na8199_9, na8200_10, na8201_9,
                   na8202_10, na8203_9, na8204_10, na8205_9, na8206_10, na8207_9, na8208_10, na8209_9, na8210_10, na8211_9, na8212_10,
                   na8213_9, na8214_10, na8215_9, na8216_10, na8217_9, na8218_10, na8219_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na8220_10, na8221_9, na8222_10, na8223_9, na8224_10, na8225_9, na8226_10, na8227_9, na8228_10, na8229_9, na8230_10,
                   na8231_9, na8232_10, na8233_9, na8234_10, na8235_9, na8236_10, na8237_9, na8238_10, na8239_9, na8240_10, na8241_9,
                   na8242_10, na8243_9, na8244_10, na8245_9, na8246_10, na8247_9, na8248_10, na8249_9, na8250_10, na8251_9, na8252_10,
                   na8253_9, na8254_10, na8255_9, na8256_10, na8257_9, na8258_10, na8259_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_///AND/      x60y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6649_4 ( .OUT(na6649_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6649_6 ( .RAM_O2(na6649_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6649_2), .COMP_OUT(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_00_16_80_B5_03_03_00_03_03_00_00_13_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6650 ( .DOA({na6650_1, na6650_2, na6650_3, na6650_4, na6650_5, na6650_6, na6650_7, na6650_8, na6650_9, na6650_10, na6650_11,
                   na6650_12, na6650_13, na6650_14, na6650_15, na6650_16, na6650_17, na6650_18, na6650_19, na6650_20, _d5045, _d5046,
                   _d5047, _d5048, _d5049, _d5050, _d5051, _d5052, _d5053, _d5054, _d5055, _d5056, na6650_33, na6650_34, na6650_35,
                   na6650_36, na6650_37, na6650_38, na6650_39, na6650_40}),
                    .DOAX({_d5057, _d5058, _d5059, _d5060, _d5061, _d5062, _d5063, _d5064, _d5065, _d5066, _d5067, _d5068, _d5069, _d5070,
                   _d5071, _d5072, _d5073, _d5074, _d5075, _d5076, _d5077, _d5078, _d5079, _d5080, _d5081, _d5082, _d5083, _d5084, _d5085,
                   _d5086, _d5087, _d5088, _d5089, _d5090, _d5091, _d5092, _d5093, _d5094, _d5095, _d5096}),
                    .DOB({_d5097, _d5098, _d5099, _d5100, _d5101, _d5102, _d5103, _d5104, _d5105, _d5106, _d5107, _d5108, _d5109, _d5110,
                   _d5111, _d5112, _d5113, _d5114, _d5115, _d5116, _d5117, _d5118, _d5119, _d5120, _d5121, _d5122, _d5123, _d5124, _d5125,
                   _d5126, _d5127, _d5128, _d5129, _d5130, _d5131, _d5132, _d5133, _d5134, _d5135, _d5136}),
                    .DOBX({_d5137, _d5138, _d5139, _d5140, _d5141, _d5142, _d5143, _d5144, _d5145, _d5146, _d5147, _d5148, _d5149, _d5150,
                   _d5151, _d5152, _d5153, _d5154, _d5155, _d5156, _d5157, _d5158, _d5159, _d5160, _d5161, _d5162, _d5163, _d5164, _d5165,
                   _d5166, _d5167, _d5168, _d5169, _d5170, _d5171, _d5172, _d5173, _d5174, _d5175, _d5176}),
                    .ECC1B_ERRA({_d5177, _d5178, _d5179, _d5180}),
                    .ECC1B_ERRB({_d5181, _d5182, _d5183, _d5184}),
                    .ECC2B_ERRA({_d5185, _d5186, _d5187, _d5188}),
                    .ECC2B_ERRB({_d5189, _d5190, _d5191, _d5192}),
                    .FORW_CAS_WRAO(_d5193), .FORW_CAS_WRBO(_d5194), .FORW_CAS_BMAO(_d5195), .FORW_CAS_BMBO(_d5196), .FORW_CAS_RDAO(_d5197),
                    .FORW_CAS_RDBO(_d5198), .FORW_UADDRAO({_d5199, _d5200, _d5201, _d5202, _d5203, _d5204, _d5205, _d5206, _d5207, _d5208,
                   _d5209, _d5210, _d5211, _d5212, _d5213, _d5214}),
                    .FORW_LADDRAO({_d5215, _d5216, _d5217, _d5218, _d5219, _d5220, _d5221, _d5222, _d5223, _d5224, _d5225, _d5226, _d5227,
                   _d5228, _d5229, _d5230}),
                    .FORW_UADDRBO({_d5231, _d5232, _d5233, _d5234, _d5235, _d5236, _d5237, _d5238, _d5239, _d5240, _d5241, _d5242, _d5243,
                   _d5244, _d5245, _d5246}),
                    .FORW_LADDRBO({_d5247, _d5248, _d5249, _d5250, _d5251, _d5252, _d5253, _d5254, _d5255, _d5256, _d5257, _d5258, _d5259,
                   _d5260, _d5261, _d5262}),
                    .FORW_UA0CLKO(_d5263), .FORW_UA0ENO(_d5264), .FORW_UA0WEO(_d5265), .FORW_LA0CLKO(_d5266), .FORW_LA0ENO(_d5267),
                    .FORW_LA0WEO(_d5268), .FORW_UA1CLKO(_d5269), .FORW_UA1ENO(_d5270), .FORW_UA1WEO(_d5271), .FORW_LA1CLKO(_d5272),
                    .FORW_LA1ENO(_d5273), .FORW_LA1WEO(_d5274), .FORW_UB0CLKO(_d5275), .FORW_UB0ENO(_d5276), .FORW_UB0WEO(_d5277), .FORW_LB0CLKO(_d5278),
                    .FORW_LB0ENO(_d5279), .FORW_LB0WEO(_d5280), .FORW_UB1CLKO(_d5281), .FORW_UB1ENO(_d5282), .FORW_UB1WEO(_d5283), .FORW_LB1CLKO(_d5284),
                    .FORW_LB1ENO(_d5285), .FORW_LB1WEO(_d5286), .CLOCKA({_d5287, _d5288, _d5289, _d5290}),
                    .CLOCKB({_d5291, _d5292, _d5293, _d5294}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, na8260_9, 1'b1, na8261_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na8262_10, 1'b1, na8263_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na8264_10, na8265_9, na8266_10, na8268_9, na8269_10, na8270_9, na8273_10, na8276_9, na8279_10, na8281_9,
                   na8282_10, na8284_9, na8290_10, na8291_9, na8293_10, na8298_9}),
                    .ADDRA1({na8299_10, na8301_9, na8303_10, na8306_9, na8308_10, na8311_9, na8316_10, na8320_9, na8321_10, na8326_9,
                   na8331_10, na8334_9, na8335_10, na8336_9, na8340_10, na8342_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8343_9, 1'b1, na8347_9, na8350_10, na8351_9, na8353_10,
                   na8354_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8356_9, 1'b1, na8359_9, na8364_10, na8366_9, na8368_10,
                   na8369_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na8374_10, na8376_9, na8380_10, na8381_9, na8497_10, na8498_9, na8499_10, na8500_9, na8501_10, na8502_9, na8503_10,
                   na8504_9, na8505_10, na8506_9, na8507_10, na8508_9, na8509_10, na8510_9, na8511_10, na8512_9, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8513_10, na8514_9, na8515_10, na8516_9, na8517_10, na8518_9, na8519_10,
                   na8520_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na8521_10, na8522_9, na8523_10, na8524_9, na8525_10, na8526_9, na8527_10, na8528_9, na8529_10, na8530_9, na8531_10,
                   na8532_9, na8533_10, na8534_9, na8535_10, na8536_9, na8537_10, na8538_9, na8539_10, na8540_9, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_00_16_80_B5_03_03_00_03_03_00_00_13_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6651 ( .DOA({na6651_1, na6651_2, na6651_3, na6651_4, na6651_5, na6651_6, na6651_7, na6651_8, na6651_9, na6651_10, na6651_11,
                   na6651_12, na6651_13, na6651_14, na6651_15, na6651_16, na6651_17, na6651_18, na6651_19, na6651_20, na6651_21, na6651_22,
                   na6651_23, na6651_24, na6651_25, na6651_26, na6651_27, na6651_28, na6651_29, na6651_30, na6651_31, na6651_32, na6651_33,
                   na6651_34, na6651_35, na6651_36, na6651_37, na6651_38, na6651_39, na6651_40}),
                    .DOAX({_d5295, _d5296, _d5297, _d5298, _d5299, _d5300, _d5301, _d5302, _d5303, _d5304, _d5305, _d5306, _d5307, _d5308,
                   _d5309, _d5310, _d5311, _d5312, _d5313, _d5314, _d5315, _d5316, _d5317, _d5318, _d5319, _d5320, _d5321, _d5322, _d5323,
                   _d5324, _d5325, _d5326, _d5327, _d5328, _d5329, _d5330, _d5331, _d5332, _d5333, _d5334}),
                    .DOB({_d5335, _d5336, _d5337, _d5338, _d5339, _d5340, _d5341, _d5342, _d5343, _d5344, _d5345, _d5346, _d5347, _d5348,
                   _d5349, _d5350, _d5351, _d5352, _d5353, _d5354, _d5355, _d5356, _d5357, _d5358, _d5359, _d5360, _d5361, _d5362, _d5363,
                   _d5364, _d5365, _d5366, _d5367, _d5368, _d5369, _d5370, _d5371, _d5372, _d5373, _d5374}),
                    .DOBX({_d5375, _d5376, _d5377, _d5378, _d5379, _d5380, _d5381, _d5382, _d5383, _d5384, _d5385, _d5386, _d5387, _d5388,
                   _d5389, _d5390, _d5391, _d5392, _d5393, _d5394, _d5395, _d5396, _d5397, _d5398, _d5399, _d5400, _d5401, _d5402, _d5403,
                   _d5404, _d5405, _d5406, _d5407, _d5408, _d5409, _d5410, _d5411, _d5412, _d5413, _d5414}),
                    .ECC1B_ERRA({_d5415, _d5416, _d5417, _d5418}),
                    .ECC1B_ERRB({_d5419, _d5420, _d5421, _d5422}),
                    .ECC2B_ERRA({_d5423, _d5424, _d5425, _d5426}),
                    .ECC2B_ERRB({_d5427, _d5428, _d5429, _d5430}),
                    .FORW_CAS_WRAO(_d5431), .FORW_CAS_WRBO(_d5432), .FORW_CAS_BMAO(_d5433), .FORW_CAS_BMBO(_d5434), .FORW_CAS_RDAO(_d5435),
                    .FORW_CAS_RDBO(_d5436), .FORW_UADDRAO({_d5437, _d5438, _d5439, _d5440, _d5441, _d5442, _d5443, _d5444, _d5445, _d5446,
                   _d5447, _d5448, _d5449, _d5450, _d5451, _d5452}),
                    .FORW_LADDRAO({_d5453, _d5454, _d5455, _d5456, _d5457, _d5458, _d5459, _d5460, _d5461, _d5462, _d5463, _d5464, _d5465,
                   _d5466, _d5467, _d5468}),
                    .FORW_UADDRBO({_d5469, _d5470, _d5471, _d5472, _d5473, _d5474, _d5475, _d5476, _d5477, _d5478, _d5479, _d5480, _d5481,
                   _d5482, _d5483, _d5484}),
                    .FORW_LADDRBO({_d5485, _d5486, _d5487, _d5488, _d5489, _d5490, _d5491, _d5492, _d5493, _d5494, _d5495, _d5496, _d5497,
                   _d5498, _d5499, _d5500}),
                    .FORW_UA0CLKO(_d5501), .FORW_UA0ENO(_d5502), .FORW_UA0WEO(_d5503), .FORW_LA0CLKO(_d5504), .FORW_LA0ENO(_d5505),
                    .FORW_LA0WEO(_d5506), .FORW_UA1CLKO(_d5507), .FORW_UA1ENO(_d5508), .FORW_UA1WEO(_d5509), .FORW_LA1CLKO(_d5510),
                    .FORW_LA1ENO(_d5511), .FORW_LA1WEO(_d5512), .FORW_UB0CLKO(_d5513), .FORW_UB0ENO(_d5514), .FORW_UB0WEO(_d5515), .FORW_LB0CLKO(_d5516),
                    .FORW_LB0ENO(_d5517), .FORW_LB0WEO(_d5518), .FORW_UB1CLKO(_d5519), .FORW_UB1ENO(_d5520), .FORW_UB1WEO(_d5521), .FORW_LB1CLKO(_d5522),
                    .FORW_LB1ENO(_d5523), .FORW_LB1WEO(_d5524), .CLOCKA({_d5525, _d5526, _d5527, _d5528}),
                    .CLOCKB({_d5529, _d5530, _d5531, _d5532}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, na8541_9, 1'b1, na8542_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na8543_10, 1'b1, na8544_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na8545_10, na8546_9, na8547_10, na8548_9, na8549_10, na8550_9, na8551_10, na8552_9, na8553_10, na8554_9,
                   na8555_10, na8556_9, na8557_10, na8558_9, na8559_10, na8560_9}),
                    .ADDRA1({na8561_10, na8562_9, na8563_10, na8564_9, na8565_10, na8566_9, na8567_10, na8568_9, na8569_10, na8570_9,
                   na8571_10, na8572_9, na8573_10, na8574_9, na8575_10, na8576_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8577_9, 1'b1, na8578_9, na8579_10, na8580_9, na8581_10,
                   na8582_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8583_9, 1'b1, na8584_9, na8585_10, na8586_9, na8587_10,
                   na8588_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na8589_10, na8590_9, na8591_10, na8592_9, na8593_10, na8594_9, na8595_10, na8596_9, na8597_10, na8598_9, na8599_10,
                   na8600_9, na8601_10, na8602_9, na8603_10, na8604_9, na8605_10, na8606_9, na8607_10, na8608_9, na8609_10, na8610_9,
                   na8611_10, na8612_9, na8613_10, na8614_9, na8615_10, na8616_9, na8617_10, na8618_9, na8619_10, na8620_9, na8621_10,
                   na8622_9, na8623_10, na8624_9, na8625_10, na8626_9, na8627_10, na8628_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na8629_10, na8630_9, na8631_10, na8632_9, na8633_10, na8634_9, na8635_10, na8636_9, na8637_10, na8638_9, na8639_10,
                   na8640_9, na8641_10, na8642_9, na8643_10, na8644_9, na8645_10, na8646_9, na8647_10, na8648_9, na8649_10, na8650_9,
                   na8651_10, na8652_9, na8653_10, na8654_9, na8655_10, na8656_9, na8657_10, na8658_9, na8659_10, na8660_9, na8661_10,
                   na8662_9, na8663_10, na8664_9, na8665_10, na8666_9, na8667_10, na8668_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_AND////      x60y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6652_1 ( .OUT(na6652_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6652_6 ( .RAM_O1(na6652_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6652_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_00_16_80_B5_03_03_00_03_03_00_00_13_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6653 ( .DOA({na6653_1, na6653_2, na6653_3, na6653_4, na6653_5, na6653_6, na6653_7, na6653_8, na6653_9, na6653_10, na6653_11,
                   na6653_12, na6653_13, na6653_14, na6653_15, na6653_16, na6653_17, na6653_18, na6653_19, na6653_20, na6653_21, na6653_22,
                   na6653_23, na6653_24, na6653_25, na6653_26, na6653_27, na6653_28, na6653_29, na6653_30, na6653_31, na6653_32, na6653_33,
                   na6653_34, na6653_35, na6653_36, na6653_37, na6653_38, na6653_39, na6653_40}),
                    .DOAX({_d5533, _d5534, _d5535, _d5536, _d5537, _d5538, _d5539, _d5540, _d5541, _d5542, _d5543, _d5544, _d5545, _d5546,
                   _d5547, _d5548, _d5549, _d5550, _d5551, _d5552, _d5553, _d5554, _d5555, _d5556, _d5557, _d5558, _d5559, _d5560, _d5561,
                   _d5562, _d5563, _d5564, _d5565, _d5566, _d5567, _d5568, _d5569, _d5570, _d5571, _d5572}),
                    .DOB({_d5573, _d5574, _d5575, _d5576, _d5577, _d5578, _d5579, _d5580, _d5581, _d5582, _d5583, _d5584, _d5585, _d5586,
                   _d5587, _d5588, _d5589, _d5590, _d5591, _d5592, _d5593, _d5594, _d5595, _d5596, _d5597, _d5598, _d5599, _d5600, _d5601,
                   _d5602, _d5603, _d5604, _d5605, _d5606, _d5607, _d5608, _d5609, _d5610, _d5611, _d5612}),
                    .DOBX({_d5613, _d5614, _d5615, _d5616, _d5617, _d5618, _d5619, _d5620, _d5621, _d5622, _d5623, _d5624, _d5625, _d5626,
                   _d5627, _d5628, _d5629, _d5630, _d5631, _d5632, _d5633, _d5634, _d5635, _d5636, _d5637, _d5638, _d5639, _d5640, _d5641,
                   _d5642, _d5643, _d5644, _d5645, _d5646, _d5647, _d5648, _d5649, _d5650, _d5651, _d5652}),
                    .ECC1B_ERRA({_d5653, _d5654, _d5655, _d5656}),
                    .ECC1B_ERRB({_d5657, _d5658, _d5659, _d5660}),
                    .ECC2B_ERRA({_d5661, _d5662, _d5663, _d5664}),
                    .ECC2B_ERRB({_d5665, _d5666, _d5667, _d5668}),
                    .FORW_CAS_WRAO(_d5669), .FORW_CAS_WRBO(_d5670), .FORW_CAS_BMAO(_d5671), .FORW_CAS_BMBO(_d5672), .FORW_CAS_RDAO(_d5673),
                    .FORW_CAS_RDBO(_d5674), .FORW_UADDRAO({_d5675, _d5676, _d5677, _d5678, _d5679, _d5680, _d5681, _d5682, _d5683, _d5684,
                   _d5685, _d5686, _d5687, _d5688, _d5689, _d5690}),
                    .FORW_LADDRAO({_d5691, _d5692, _d5693, _d5694, _d5695, _d5696, _d5697, _d5698, _d5699, _d5700, _d5701, _d5702, _d5703,
                   _d5704, _d5705, _d5706}),
                    .FORW_UADDRBO({_d5707, _d5708, _d5709, _d5710, _d5711, _d5712, _d5713, _d5714, _d5715, _d5716, _d5717, _d5718, _d5719,
                   _d5720, _d5721, _d5722}),
                    .FORW_LADDRBO({_d5723, _d5724, _d5725, _d5726, _d5727, _d5728, _d5729, _d5730, _d5731, _d5732, _d5733, _d5734, _d5735,
                   _d5736, _d5737, _d5738}),
                    .FORW_UA0CLKO(_d5739), .FORW_UA0ENO(_d5740), .FORW_UA0WEO(_d5741), .FORW_LA0CLKO(_d5742), .FORW_LA0ENO(_d5743),
                    .FORW_LA0WEO(_d5744), .FORW_UA1CLKO(_d5745), .FORW_UA1ENO(_d5746), .FORW_UA1WEO(_d5747), .FORW_LA1CLKO(_d5748),
                    .FORW_LA1ENO(_d5749), .FORW_LA1WEO(_d5750), .FORW_UB0CLKO(_d5751), .FORW_UB0ENO(_d5752), .FORW_UB0WEO(_d5753), .FORW_LB0CLKO(_d5754),
                    .FORW_LB0ENO(_d5755), .FORW_LB0WEO(_d5756), .FORW_UB1CLKO(_d5757), .FORW_UB1ENO(_d5758), .FORW_UB1WEO(_d5759), .FORW_LB1CLKO(_d5760),
                    .FORW_LB1ENO(_d5761), .FORW_LB1WEO(_d5762), .CLOCKA({_d5763, _d5764, _d5765, _d5766}),
                    .CLOCKB({_d5767, _d5768, _d5769, _d5770}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, na8669_9, 1'b1, na8670_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na8671_10, 1'b1, na8672_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na8673_10, na8674_9, na8675_10, na8676_9, na8677_10, na8678_9, na8679_10, na8680_9, na8681_10, na8682_9,
                   na8683_10, na8684_9, na8685_10, na8686_9, na8687_10, na8688_9}),
                    .ADDRA1({na8689_10, na8690_9, na8691_10, na8692_9, na8693_10, na8694_9, na8695_10, na8696_9, na8697_10, na8698_9,
                   na8699_10, na8700_9, na8701_10, na8702_9, na8703_10, na8704_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8705_9, 1'b1, na8706_9, na8707_10, na8708_9, na8709_10,
                   na8710_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8711_9, 1'b1, na8712_9, na8713_10, na8714_9, na8715_10,
                   na8716_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na8717_10, na8718_9, na8719_10, na8720_9, na8721_10, na8722_9, na8723_10, na8724_9, na8725_10, na8726_9, na8727_10,
                   na8728_9, na8729_10, na8730_9, na8731_10, na8732_9, na8733_10, na8734_9, na8735_10, na8736_9, na8737_10, na8738_9,
                   na8739_10, na8740_9, na8741_10, na8742_9, na8743_10, na8744_9, na8745_10, na8746_9, na8747_10, na8748_9, na8749_10,
                   na8750_9, na8751_10, na8752_9, na8753_10, na8754_9, na8755_10, na8756_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na8757_10, na8758_9, na8759_10, na8760_9, na8761_10, na8762_9, na8763_10, na8764_9, na8765_10, na8766_9, na8767_10,
                   na8768_9, na8769_10, na8770_9, na8771_10, na8772_9, na8773_10, na8774_9, na8775_10, na8776_9, na8777_10, na8778_9,
                   na8779_10, na8780_9, na8781_10, na8782_9, na8783_10, na8784_9, na8785_10, na8786_9, na8787_10, na8788_9, na8789_10,
                   na8790_9, na8791_10, na8792_9, na8793_10, na8794_9, na8795_10, na8796_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_///AND/      x60y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6654_4 ( .OUT(na6654_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6654_6 ( .RAM_O2(na6654_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6654_2), .COMP_OUT(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_05_00_02_80_15_00_00_00_03_03_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6655 ( .DOA({_d5771, _d5772, _d5773, _d5774, _d5775, _d5776, _d5777, _d5778, _d5779, _d5780, _d5781, _d5782, _d5783, _d5784,
                   _d5785, _d5786, _d5787, _d5788, _d5789, _d5790, na6655_21, na6655_22, na6655_23, na6655_24, na6655_25, na6655_26,
                   na6655_27, na6655_28, na6655_29, na6655_30, na6655_31, na6655_32, na6655_33, na6655_34, na6655_35, na6655_36, na6655_37,
                   na6655_38, na6655_39, na6655_40}),
                    .DOAX({_d5791, _d5792, _d5793, _d5794, _d5795, _d5796, _d5797, _d5798, _d5799, _d5800, _d5801, _d5802, _d5803, _d5804,
                   _d5805, _d5806, _d5807, _d5808, _d5809, _d5810, _d5811, _d5812, _d5813, _d5814, _d5815, _d5816, _d5817, _d5818, _d5819,
                   _d5820, _d5821, _d5822, _d5823, _d5824, _d5825, _d5826, _d5827, _d5828, _d5829, _d5830}),
                    .DOB({_d5831, _d5832, _d5833, _d5834, _d5835, _d5836, _d5837, _d5838, _d5839, _d5840, _d5841, _d5842, _d5843, _d5844,
                   _d5845, _d5846, _d5847, _d5848, _d5849, _d5850, _d5851, _d5852, _d5853, _d5854, _d5855, _d5856, _d5857, _d5858, _d5859,
                   _d5860, _d5861, _d5862, _d5863, _d5864, _d5865, _d5866, _d5867, _d5868, _d5869, _d5870}),
                    .DOBX({_d5871, _d5872, _d5873, _d5874, _d5875, _d5876, _d5877, _d5878, _d5879, _d5880, _d5881, _d5882, _d5883, _d5884,
                   _d5885, _d5886, _d5887, _d5888, _d5889, _d5890, _d5891, _d5892, _d5893, _d5894, _d5895, _d5896, _d5897, _d5898, _d5899,
                   _d5900, _d5901, _d5902, _d5903, _d5904, _d5905, _d5906, _d5907, _d5908, _d5909, _d5910}),
                    .ECC1B_ERRA({_d5911, _d5912, _d5913, _d5914}),
                    .ECC1B_ERRB({_d5915, _d5916, _d5917, _d5918}),
                    .ECC2B_ERRA({_d5919, _d5920, _d5921, _d5922}),
                    .ECC2B_ERRB({_d5923, _d5924, _d5925, _d5926}),
                    .FORW_CAS_WRAO(_d5927), .FORW_CAS_WRBO(_d5928), .FORW_CAS_BMAO(_d5929), .FORW_CAS_BMBO(_d5930), .FORW_CAS_RDAO(_d5931),
                    .FORW_CAS_RDBO(_d5932), .FORW_UADDRAO({_d5933, _d5934, _d5935, _d5936, _d5937, _d5938, _d5939, _d5940, _d5941, _d5942,
                   _d5943, _d5944, _d5945, _d5946, _d5947, _d5948}),
                    .FORW_LADDRAO({_d5949, _d5950, _d5951, _d5952, _d5953, _d5954, _d5955, _d5956, _d5957, _d5958, _d5959, _d5960, _d5961,
                   _d5962, _d5963, _d5964}),
                    .FORW_UADDRBO({_d5965, _d5966, _d5967, _d5968, _d5969, _d5970, _d5971, _d5972, _d5973, _d5974, _d5975, _d5976, _d5977,
                   _d5978, _d5979, _d5980}),
                    .FORW_LADDRBO({_d5981, _d5982, _d5983, _d5984, _d5985, _d5986, _d5987, _d5988, _d5989, _d5990, _d5991, _d5992, _d5993,
                   _d5994, _d5995, _d5996}),
                    .FORW_UA0CLKO(_d5997), .FORW_UA0ENO(_d5998), .FORW_UA0WEO(_d5999), .FORW_LA0CLKO(_d6000), .FORW_LA0ENO(_d6001),
                    .FORW_LA0WEO(_d6002), .FORW_UA1CLKO(_d6003), .FORW_UA1ENO(_d6004), .FORW_UA1WEO(_d6005), .FORW_LA1CLKO(_d6006),
                    .FORW_LA1ENO(_d6007), .FORW_LA1WEO(_d6008), .FORW_UB0CLKO(_d6009), .FORW_UB0ENO(_d6010), .FORW_UB0WEO(_d6011), .FORW_LB0CLKO(_d6012),
                    .FORW_LB0ENO(_d6013), .FORW_LB0WEO(_d6014), .FORW_UB1CLKO(_d6015), .FORW_UB1ENO(_d6016), .FORW_UB1WEO(_d6017), .FORW_LB1CLKO(_d6018),
                    .FORW_LB1ENO(_d6019), .FORW_LB1WEO(_d6020), .CLOCKA({_d6021, _d6022, _d6023, _d6024}),
                    .CLOCKB({_d6025, _d6026, _d6027, _d6028}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, na8797_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, 1'b1, 1'b1, na8798_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na8799_10, na8800_9, na8801_10, na8802_9, na8803_10, na8804_9, na8805_10, na8806_9, na8807_10, na8808_9,
                   na8809_10, na8810_9, na8811_10, na8812_9, na8813_10, na8814_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8815_9, 1'b1, na8816_9, na8817_10, na8818_9, na8819_10,
                   na8820_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na8821_10, na8822_9, na8823_10, na8824_9, na8825_10, na8826_9, na8827_10, na8828_9, na8829_10, na8830_9,
                   na8831_10, na8832_9, na8833_10, na8834_9, na8835_10, na8836_9, na8837_10, na8838_9, na8839_10, na8840_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na8841_10, na8842_9, na8843_10, na8844_9, na8845_10, na8846_9, na8847_10, na8848_9, na8849_10, na8850_9,
                   na8851_10, na8852_9, na8853_10, na8854_9, na8855_10, na8856_9, na8857_10, na8858_9, na8859_10, na8860_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_AND////      x60y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6656_1 ( .OUT(na6656_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6656_6 ( .RAM_O1(na6656_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6656_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_00_16_80_B5_03_03_00_03_03_00_00_13_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6657 ( .DOA({na6657_1, na6657_2, na6657_3, na6657_4, na6657_5, na6657_6, na6657_7, na6657_8, na6657_9, na6657_10, na6657_11,
                   na6657_12, na6657_13, na6657_14, na6657_15, na6657_16, na6657_17, na6657_18, na6657_19, na6657_20, na6657_21, na6657_22,
                   na6657_23, na6657_24, na6657_25, na6657_26, na6657_27, na6657_28, na6657_29, na6657_30, na6657_31, na6657_32, na6657_33,
                   na6657_34, na6657_35, na6657_36, na6657_37, na6657_38, na6657_39, na6657_40}),
                    .DOAX({_d6029, _d6030, _d6031, _d6032, _d6033, _d6034, _d6035, _d6036, _d6037, _d6038, _d6039, _d6040, _d6041, _d6042,
                   _d6043, _d6044, _d6045, _d6046, _d6047, _d6048, _d6049, _d6050, _d6051, _d6052, _d6053, _d6054, _d6055, _d6056, _d6057,
                   _d6058, _d6059, _d6060, _d6061, _d6062, _d6063, _d6064, _d6065, _d6066, _d6067, _d6068}),
                    .DOB({_d6069, _d6070, _d6071, _d6072, _d6073, _d6074, _d6075, _d6076, _d6077, _d6078, _d6079, _d6080, _d6081, _d6082,
                   _d6083, _d6084, _d6085, _d6086, _d6087, _d6088, _d6089, _d6090, _d6091, _d6092, _d6093, _d6094, _d6095, _d6096, _d6097,
                   _d6098, _d6099, _d6100, _d6101, _d6102, _d6103, _d6104, _d6105, _d6106, _d6107, _d6108}),
                    .DOBX({_d6109, _d6110, _d6111, _d6112, _d6113, _d6114, _d6115, _d6116, _d6117, _d6118, _d6119, _d6120, _d6121, _d6122,
                   _d6123, _d6124, _d6125, _d6126, _d6127, _d6128, _d6129, _d6130, _d6131, _d6132, _d6133, _d6134, _d6135, _d6136, _d6137,
                   _d6138, _d6139, _d6140, _d6141, _d6142, _d6143, _d6144, _d6145, _d6146, _d6147, _d6148}),
                    .ECC1B_ERRA({_d6149, _d6150, _d6151, _d6152}),
                    .ECC1B_ERRB({_d6153, _d6154, _d6155, _d6156}),
                    .ECC2B_ERRA({_d6157, _d6158, _d6159, _d6160}),
                    .ECC2B_ERRB({_d6161, _d6162, _d6163, _d6164}),
                    .FORW_CAS_WRAO(_d6165), .FORW_CAS_WRBO(_d6166), .FORW_CAS_BMAO(_d6167), .FORW_CAS_BMBO(_d6168), .FORW_CAS_RDAO(_d6169),
                    .FORW_CAS_RDBO(_d6170), .FORW_UADDRAO({_d6171, _d6172, _d6173, _d6174, _d6175, _d6176, _d6177, _d6178, _d6179, _d6180,
                   _d6181, _d6182, _d6183, _d6184, _d6185, _d6186}),
                    .FORW_LADDRAO({_d6187, _d6188, _d6189, _d6190, _d6191, _d6192, _d6193, _d6194, _d6195, _d6196, _d6197, _d6198, _d6199,
                   _d6200, _d6201, _d6202}),
                    .FORW_UADDRBO({_d6203, _d6204, _d6205, _d6206, _d6207, _d6208, _d6209, _d6210, _d6211, _d6212, _d6213, _d6214, _d6215,
                   _d6216, _d6217, _d6218}),
                    .FORW_LADDRBO({_d6219, _d6220, _d6221, _d6222, _d6223, _d6224, _d6225, _d6226, _d6227, _d6228, _d6229, _d6230, _d6231,
                   _d6232, _d6233, _d6234}),
                    .FORW_UA0CLKO(_d6235), .FORW_UA0ENO(_d6236), .FORW_UA0WEO(_d6237), .FORW_LA0CLKO(_d6238), .FORW_LA0ENO(_d6239),
                    .FORW_LA0WEO(_d6240), .FORW_UA1CLKO(_d6241), .FORW_UA1ENO(_d6242), .FORW_UA1WEO(_d6243), .FORW_LA1CLKO(_d6244),
                    .FORW_LA1ENO(_d6245), .FORW_LA1WEO(_d6246), .FORW_UB0CLKO(_d6247), .FORW_UB0ENO(_d6248), .FORW_UB0WEO(_d6249), .FORW_LB0CLKO(_d6250),
                    .FORW_LB0ENO(_d6251), .FORW_LB0WEO(_d6252), .FORW_UB1CLKO(_d6253), .FORW_UB1ENO(_d6254), .FORW_UB1WEO(_d6255), .FORW_LB1CLKO(_d6256),
                    .FORW_LB1ENO(_d6257), .FORW_LB1WEO(_d6258), .CLOCKA({_d6259, _d6260, _d6261, _d6262}),
                    .CLOCKB({_d6263, _d6264, _d6265, _d6266}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, na8861_9, 1'b1, na8862_9}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na8863_10, 1'b1, na8864_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na8865_10, na8866_9, na8867_10, na8868_9, na8869_10, na8870_9, na8871_10, na8872_9, na8873_10, na8874_9,
                   na8875_10, na8876_9, na8877_10, na8878_9, na8879_10, na8880_9}),
                    .ADDRA1({na8881_10, na8882_9, na8883_10, na8884_9, na8885_10, na8886_9, na8887_10, na8888_9, na8889_10, na8890_9,
                   na8891_10, na8892_9, na8893_10, na8894_9, na8895_10, na8896_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8897_9, 1'b1, na8898_9, na8899_10, na8900_9, na8901_10,
                   na8902_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na8903_9, 1'b1, na8904_9, na8905_10, na8906_9, na8907_10,
                   na8908_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na8909_10, na8910_9, na8911_10, na8912_9, na8913_10, na8914_9, na8915_10, na8916_9, na8917_10, na8918_9, na8919_10,
                   na8920_9, na8921_10, na8922_9, na8923_10, na8924_9, na8925_10, na8926_9, na8927_10, na8928_9, na8929_10, na8930_9,
                   na8931_10, na8932_9, na8933_10, na8934_9, na8935_10, na8936_9, na8937_10, na8938_9, na8939_10, na8940_9, na8941_10,
                   na8942_9, na8943_10, na8944_9, na8945_10, na8946_9, na8947_10, na8948_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na8949_10, na8950_9, na8951_10, na8952_9, na8953_10, na8954_9, na8955_10, na8956_9, na8957_10, na8958_9, na8959_10,
                   na8960_9, na8961_10, na8962_9, na8963_10, na8964_9, na8965_10, na8966_9, na8967_10, na8968_9, na8969_10, na8970_9,
                   na8971_10, na8972_9, na8973_10, na8974_9, na8975_10, na8976_9, na8977_10, na8978_9, na8979_10, na8980_9, na8981_10,
                   na8982_9, na8983_10, na8984_9, na8985_10, na8986_9, na8987_10, na8988_9}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_///AND/      x60y70     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6658_4 ( .OUT(na6658_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2518_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6658_6 ( .RAM_O2(na6658_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6658_2), .COMP_OUT(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_04_80_00_91_03_00_23_03_00_23_00_13_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a6659 ( .DOA({_d6267, _d6268, _d6269, _d6270, _d6271, _d6272, _d6273, _d6274, _d6275, _d6276, _d6277, _d6278, _d6279, _d6280,
                   _d6281, _d6282, _d6283, _d6284, _d6285, _d6286, _d6287, _d6288, _d6289, _d6290, _d6291, _d6292, _d6293, _d6294, _d6295,
                   _d6296, _d6297, _d6298, _d6299, _d6300, _d6301, _d6302, _d6303, _d6304, _d6305, _d6306}),
                    .DOAX({_d6307, _d6308, _d6309, _d6310, _d6311, _d6312, _d6313, _d6314, _d6315, _d6316, _d6317, _d6318, _d6319, _d6320,
                   _d6321, _d6322, _d6323, _d6324, _d6325, _d6326, _d6327, _d6328, _d6329, _d6330, _d6331, _d6332, _d6333, _d6334, _d6335,
                   _d6336, _d6337, _d6338, _d6339, _d6340, _d6341, _d6342, _d6343, _d6344, _d6345, _d6346}),
                    .DOB({_d6347, _d6348, _d6349, _d6350, _d6351, _d6352, _d6353, _d6354, _d6355, _d6356, _d6357, _d6358, na6659_93,
                   na6659_94, na6659_95, na6659_96, na6659_97, na6659_98, na6659_99, na6659_100, _d6359, _d6360, _d6361, _d6362, _d6363,
                   _d6364, _d6365, _d6366, _d6367, _d6368, _d6369, _d6370, na6659_113, na6659_114, na6659_115, na6659_116, na6659_117,
                   na6659_118, na6659_119, na6659_120}),
                    .DOBX({_d6371, _d6372, _d6373, _d6374, _d6375, _d6376, _d6377, _d6378, _d6379, _d6380, _d6381, _d6382, _d6383, _d6384,
                   _d6385, _d6386, _d6387, _d6388, _d6389, _d6390, _d6391, _d6392, _d6393, _d6394, _d6395, _d6396, _d6397, _d6398, _d6399,
                   _d6400, _d6401, _d6402, _d6403, _d6404, _d6405, _d6406, _d6407, _d6408, _d6409, _d6410}),
                    .ECC1B_ERRA({_d6411, _d6412, _d6413, _d6414}),
                    .ECC1B_ERRB({_d6415, _d6416, _d6417, _d6418}),
                    .ECC2B_ERRA({_d6419, _d6420, _d6421, _d6422}),
                    .ECC2B_ERRB({_d6423, _d6424, _d6425, _d6426}),
                    .FORW_CAS_WRAO(_d6427), .FORW_CAS_WRBO(_d6428), .FORW_CAS_BMAO(_d6429), .FORW_CAS_BMBO(_d6430), .FORW_CAS_RDAO(_d6431),
                    .FORW_CAS_RDBO(_d6432), .FORW_UADDRAO({_d6433, _d6434, _d6435, _d6436, _d6437, _d6438, _d6439, _d6440, _d6441, _d6442,
                   _d6443, _d6444, _d6445, _d6446, _d6447, _d6448}),
                    .FORW_LADDRAO({_d6449, _d6450, _d6451, _d6452, _d6453, _d6454, _d6455, _d6456, _d6457, _d6458, _d6459, _d6460, _d6461,
                   _d6462, _d6463, _d6464}),
                    .FORW_UADDRBO({_d6465, _d6466, _d6467, _d6468, _d6469, _d6470, _d6471, _d6472, _d6473, _d6474, _d6475, _d6476, _d6477,
                   _d6478, _d6479, _d6480}),
                    .FORW_LADDRBO({_d6481, _d6482, _d6483, _d6484, _d6485, _d6486, _d6487, _d6488, _d6489, _d6490, _d6491, _d6492, _d6493,
                   _d6494, _d6495, _d6496}),
                    .FORW_UA0CLKO(_d6497), .FORW_UA0ENO(_d6498), .FORW_UA0WEO(_d6499), .FORW_LA0CLKO(_d6500), .FORW_LA0ENO(_d6501),
                    .FORW_LA0WEO(_d6502), .FORW_UA1CLKO(_d6503), .FORW_UA1ENO(_d6504), .FORW_UA1WEO(_d6505), .FORW_LA1CLKO(_d6506),
                    .FORW_LA1ENO(_d6507), .FORW_LA1WEO(_d6508), .FORW_UB0CLKO(_d6509), .FORW_UB0ENO(_d6510), .FORW_UB0WEO(_d6511), .FORW_LB0CLKO(_d6512),
                    .FORW_LB0ENO(_d6513), .FORW_LB0WEO(_d6514), .FORW_UB1CLKO(_d6515), .FORW_UB1ENO(_d6516), .FORW_UB1WEO(_d6517), .FORW_LB1CLKO(_d6518),
                    .FORW_LB1ENO(_d6519), .FORW_LB1WEO(_d6520), .CLOCKA({_d6521, _d6522, _d6523, _d6524}),
                    .CLOCKB({_d6525, _d6526, _d6527, _d6528}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, na8989_9, 1'b1, na8990_9}),
                    .GLWEA({1'b1, na8991_10, 1'b1, na8992_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na8993_10, na8994_9, na8995_10, na8996_9, na8997_10, na8998_9, na8999_10, na9000_9, na9001_10, na9002_9,
                   na9003_10, na9004_9, na9005_10, na9006_9, na9007_10, na9008_9}),
                    .ADDRA1({na9009_10, na9010_9, na9011_10, na9012_9, na9013_10, na9014_9, na9015_10, na9016_9, na9017_10, na9018_9,
                   na9019_10, na9020_9, na9021_10, na9022_9, na9023_10, na9024_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({na9025_10, na9026_9, na9027_10, na9028_9, na9029_10, na9030_9, na9031_10, na9032_9, na9033_10, na9034_9,
                   na9035_10, na9036_9, na9037_10, na9038_9, na9039_10, na9040_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({na9041_10, na9042_9, na9043_10, na9044_9, na9045_10, na9046_9, na9047_10, na9048_9, na9049_10, na9050_9,
                   na9051_10, na9052_9, na9053_10, na9054_9, na9055_10, na9056_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na9057_10, na9058_9, na9059_10, na9060_9, na9061_10, na9062_9, na9063_10, na9064_9, na9065_10, na9066_9, na9067_10,
                   na9068_9, na9069_10, na9070_9, na9071_10, na9072_9, na9073_10, na9074_9, na9075_10, na9076_9, na9077_10, na9078_9,
                   na9079_10, na9080_9, na9081_10, na9082_9, na9083_10, na9084_9, na9085_10, na9086_9, na9087_10, na9088_9, na9089_10,
                   na9090_9, na9091_10, na9092_9, na9093_10, na9094_9, na9095_10, na9096_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na9097_10, na9098_9, na9099_10, na9100_9, na9101_10, na9102_9, na9103_10, na9104_9, na9105_10, na9106_9, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na9107_10, na9108_9, na9109_10, na9110_9, na9111_10, na9112_9,
                   na9113_10, na9114_9, na9115_10, na9116_9, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na4116_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_AND////      x60y70     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6660_1 ( .OUT(na6660_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2517_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6660_6 ( .RAM_O1(na6660_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6660_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_////RAM_I2      x1y128     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6661_5 ( .OUT(na6661_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6627_2), .CP_O(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a6662 ( .PCLK0(na6662_1), .PCLK1(_d6529), .PCLK2(_d6530), .PCLK3(_d6531), .CLK0(na6570_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                    .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_AND////      x68y80     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6663_1 ( .OUT(na6663_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9827_2), .IN6(1'b1), .IN7(na517_2), .IN8(na3950_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x49y69     80'h00_0018_00_0000_0EEE_0757
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6664_1 ( .OUT(na6664_1), .IN1(~na3487_1), .IN2(~na9152_2), .IN3(~na3491_1), .IN4(1'b0), .IN5(~na50_1), .IN6(~na3489_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x1y66     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6665_5 ( .OUT(na6665_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6628_1), .CP_O(1'b0) );
// C_///OR/      x51y50     80'h00_0060_00_0000_0C0E_FF5B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a6666_4 ( .OUT(na6666_2), .IN1(na9207_2), .IN2(~na5948_1), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y69     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6667_4 ( .OUT(na6667_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2516_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6667_6 ( .RAM_O2(na6667_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6667_2), .COMP_OUT(1'b0) );
// C_OR////      x50y52     80'h00_0018_00_0000_0CEE_7C00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6668_1 ( .OUT(na6668_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na369_2), .IN7(~na3268_2), .IN8(~na5962_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y69     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6669_1 ( .OUT(na6669_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2515_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6669_6 ( .RAM_O1(na6669_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6669_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y68     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6670_4 ( .OUT(na6670_2), .IN1(na2514_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6670_6 ( .RAM_O2(na6670_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6670_2), .COMP_OUT(1'b0) );
// C_///XOR/      x50y87     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6671_4 ( .OUT(na6671_2), .IN1(na3326_2), .IN2(1'b0), .IN3(na3266_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y53     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6672_1 ( .OUT(na6672_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2991_1), .IN6(1'b1), .IN7(1'b1), .IN8(na9125_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x114y40     80'h00_0078_00_0000_0C88_F4C8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6673_1 ( .OUT(na6673_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9947_2), .IN6(na36_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6673_4 ( .OUT(na6673_2), .IN1(na9_1), .IN2(na31_2), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x98y72     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6674_4 ( .OUT(na6674_2), .IN1(na9947_2), .IN2(~na36_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y65     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6675_4 ( .OUT(na6675_2), .IN1(na9947_2), .IN2(na36_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6676_1 ( .OUT(na6676_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6676_6 ( .RAM_O1(na6676_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6676_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y68     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6677_4 ( .OUT(na6677_2), .IN1(~na9947_2), .IN2(~na36_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y70     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6678_1 ( .OUT(na6678_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9947_2), .IN6(na36_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y67     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6679_4 ( .OUT(na6679_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6679_6 ( .RAM_O2(na6679_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6679_2), .COMP_OUT(1'b0) );
// C_AND////      x60y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6680_1 ( .OUT(na6680_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6680_6 ( .RAM_O1(na6680_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6680_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x103y64     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6681_1 ( .OUT(na6681_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na9947_2), .IN6(~na36_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6682_4 ( .OUT(na6682_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6682_6 ( .RAM_O2(na6682_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6682_2), .COMP_OUT(1'b0) );
// C_AND////      x60y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6683_1 ( .OUT(na6683_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6683_6 ( .RAM_O1(na6683_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6683_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x108y43     80'h00_0078_00_0000_0C88_33A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6684_1 ( .OUT(na6684_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na36_1), .IN7(1'b1), .IN8(~na6673_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6684_4 ( .OUT(na6684_2), .IN1(na9_1), .IN2(na31_2), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6685_4 ( .OUT(na6685_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6685_6 ( .RAM_O2(na6685_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6685_2), .COMP_OUT(1'b0) );
// C_AND////      x60y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6686_1 ( .OUT(na6686_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6686_6 ( .RAM_O1(na6686_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6686_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6687_4 ( .OUT(na6687_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6687_6 ( .RAM_O2(na6687_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6687_2), .COMP_OUT(1'b0) );
// C_AND////      x69y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6688_1 ( .OUT(na6688_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6688_6 ( .RAM_O1(na6688_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6688_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6689_4 ( .OUT(na6689_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6689_6 ( .RAM_O2(na6689_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6689_2), .COMP_OUT(1'b0) );
// C_AND////      x69y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6690_1 ( .OUT(na6690_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6690_6 ( .RAM_O1(na6690_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6690_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y70     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6691_4 ( .OUT(na6691_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2592_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6691_6 ( .RAM_O2(na6691_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6691_2), .COMP_OUT(1'b0) );
// C_MX2b////      x90y86     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6692_1 ( .OUT(na6692_1), .IN1(1'b1), .IN2(na2935_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1002_1), .IN8(~na2979_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y70     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6693_1 ( .OUT(na6693_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2590_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6693_6 ( .RAM_O1(na6693_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6693_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y69     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6694_4 ( .OUT(na6694_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2588_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6694_6 ( .RAM_O2(na6694_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6694_2), .COMP_OUT(1'b0) );
// C_ORAND////      x97y96     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6695_1 ( .OUT(na6695_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na114_1), .IN7(~na2937_2), .IN8(na6702_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x104y72     80'h00_0018_00_0000_0EEE_5E5A
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6696_1 ( .OUT(na6696_1), .IN1(na6699_2), .IN2(1'b0), .IN3(~na6700_2), .IN4(1'b0), .IN5(na112_2), .IN6(na6701_2), .IN7(~na6700_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y69     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6697_1 ( .OUT(na6697_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2586_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6697_6 ( .RAM_O1(na6697_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6697_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y68     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6698_4 ( .OUT(na6698_2), .IN1(na2584_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6698_6 ( .RAM_O2(na6698_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6698_2), .COMP_OUT(1'b0) );
// C_///AND/      x85y73     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6699_4 ( .OUT(na6699_2), .IN1(na95_2), .IN2(na89_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y79     80'h00_0078_00_0000_0CEE_70D0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6700_1 ( .OUT(na6700_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na97_1), .IN8(~na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a6700_4 ( .OUT(na6700_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na97_2), .IN4(na28_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y72     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6701_4 ( .OUT(na6701_2), .IN1(1'b1), .IN2(na9153_2), .IN3(1'b1), .IN4(na101_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y88     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6702_1 ( .OUT(na6702_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2978_1), .IN8(~na1001_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6703_1 ( .OUT(na6703_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6703_6 ( .RAM_O1(na6703_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6703_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y67     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6704_4 ( .OUT(na6704_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6704_6 ( .RAM_O2(na6704_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6704_2), .COMP_OUT(1'b0) );
// C_ORAND////      x95y98     80'h00_0018_00_0000_0C88_DAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6705_1 ( .OUT(na6705_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na122_1), .IN6(1'b0), .IN7(~na2937_2), .IN8(na6712_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x78y84     80'h00_0018_00_0000_0EEE_A3CB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6706_1 ( .OUT(na6706_1), .IN1(na6709_1), .IN2(~na6710_2), .IN3(1'b0), .IN4(na120_2), .IN5(1'b0), .IN6(~na6710_1), .IN7(na6711_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6707_1 ( .OUT(na6707_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6707_6 ( .RAM_O1(na6707_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6707_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6708_4 ( .OUT(na6708_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6708_6 ( .RAM_O2(na6708_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6708_2), .COMP_OUT(1'b0) );
// C_AND////      x87y79     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6709_1 ( .OUT(na6709_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na95_2), .IN6(1'b1), .IN7(na90_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x85y82     80'h00_0078_00_0000_0CEE_535A
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6710_1 ( .OUT(na6710_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na35_1), .IN7(~na97_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a6710_4 ( .OUT(na6710_2), .IN1(na29_1), .IN2(1'b0), .IN3(~na97_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y69     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6711_1 ( .OUT(na6711_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(na101_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y90     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6712_1 ( .OUT(na6712_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na9728_2), .IN8(~na1000_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6713_1 ( .OUT(na6713_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6713_6 ( .RAM_O1(na6713_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6713_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6714_4 ( .OUT(na6714_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6714_6 ( .RAM_O2(na6714_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6714_2), .COMP_OUT(1'b0) );
// C_AND////      x69y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6715_1 ( .OUT(na6715_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6715_6 ( .RAM_O1(na6715_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6715_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y72     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6716_4 ( .OUT(na6716_2_i), .IN1(na2488_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6716_5 ( .OUT(na6716_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6716_6 ( .RAM_O2(na6716_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6716_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y72     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6717_1 ( .OUT(na6717_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2486_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6717_2 ( .OUT(na6717_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6717_6 ( .RAM_O1(na6717_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6717_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y71     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6718_4 ( .OUT(na6718_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2484_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6718_5 ( .OUT(na6718_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6718_6 ( .RAM_O2(na6718_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6718_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x83y82     80'h00_0018_00_0000_0888_FD7D
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6719_1 ( .OUT(na6719_1), .IN1(~na95_2), .IN2(na9137_2), .IN3(~na84_1), .IN4(~na9175_2), .IN5(~na95_1), .IN6(na24_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x62y71     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6720_1 ( .OUT(na6720_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2480_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6720_2 ( .OUT(na6720_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6720_6 ( .RAM_O1(na6720_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6720_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y72     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6721_4 ( .OUT(na6721_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2477_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6721_5 ( .OUT(na6721_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6721_6 ( .RAM_O2(na6721_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6721_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y72     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6722_1 ( .OUT(na6722_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2474_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6722_2 ( .OUT(na6722_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6722_6 ( .RAM_O1(na6722_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6722_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x93y96     80'h00_0018_00_0000_0C88_DAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6723_1 ( .OUT(na6723_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na133_1), .IN6(1'b0), .IN7(~na2937_2), .IN8(na6724_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y86     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6724_1 ( .OUT(na6724_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2975_1), .IN6(~na2969_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y71     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6725_4 ( .OUT(na6725_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2471_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6725_5 ( .OUT(na6725_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6725_6 ( .RAM_O2(na6725_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6725_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y71     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6726_1 ( .OUT(na6726_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2468_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6726_2 ( .OUT(na6726_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6726_6 ( .RAM_O1(na6726_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6726_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND///ORAND/      x102y88     80'h00_0078_00_0000_0C88_DA5B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6727_1 ( .OUT(na6727_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na140_1), .IN6(1'b0), .IN7(~na2937_2), .IN8(na6733_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a6727_4 ( .OUT(na6727_2), .IN1(na138_1), .IN2(~na99_2), .IN3(~na97_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y70     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6728_4 ( .OUT(na6728_2_i), .IN1(1'b1), .IN2(na2465_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6728_5 ( .OUT(na6728_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6728_6 ( .RAM_O2(na6728_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6728_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y70     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6729_1 ( .OUT(na6729_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2462_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6729_2 ( .OUT(na6729_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6729_6 ( .RAM_O1(na6729_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6729_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y69     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6730_4 ( .OUT(na6730_2_i), .IN1(1'b1), .IN2(na2459_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6730_5 ( .OUT(na6730_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6730_6 ( .RAM_O2(na6730_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6730_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y69     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6731_1 ( .OUT(na6731_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2455_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6731_2 ( .OUT(na6731_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6731_6 ( .RAM_O1(na6731_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6731_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y68     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6732_4 ( .OUT(na6732_2_i), .IN1(1'b1), .IN2(na2454_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6732_5 ( .OUT(na6732_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6732_6 ( .RAM_O2(na6732_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6732_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x90y82     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6733_1 ( .OUT(na6733_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na9714_2), .IN5(1'b0), .IN6(~na962_1), .IN7(1'b0), .IN8(~na2974_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y68     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6734_1 ( .OUT(na6734_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3583_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6734_2 ( .OUT(na6734_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6734_6 ( .RAM_O1(na6734_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6734_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y67     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6735_4 ( .OUT(na6735_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3580_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6735_5 ( .OUT(na6735_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6735_6 ( .RAM_O2(na6735_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6735_2_i), .COMP_OUT(1'b0) );
// C_///ORAND/      x93y92     80'h00_0060_00_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a6736_4 ( .OUT(na6736_2), .IN1(1'b0), .IN2(na147_1), .IN3(~na2937_2), .IN4(na6741_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y67     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6737_1 ( .OUT(na6737_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3577_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6737_2 ( .OUT(na6737_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6737_6 ( .RAM_O1(na6737_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6737_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y66     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6738_4 ( .OUT(na6738_2_i), .IN1(1'b1), .IN2(na3574_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6738_5 ( .OUT(na6738_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6738_6 ( .RAM_O2(na6738_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6738_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y66     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6739_1 ( .OUT(na6739_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3571_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6739_2 ( .OUT(na6739_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6739_6 ( .RAM_O1(na6739_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6739_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y65     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6740_4 ( .OUT(na6740_2_i), .IN1(na3568_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6740_5 ( .OUT(na6740_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6740_6 ( .RAM_O2(na6740_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6740_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x94y86     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6741_1 ( .OUT(na6741_1), .IN1(1'b1), .IN2(~na2935_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1085_1), .IN8(~na921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y65     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6742_1 ( .OUT(na6742_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3565_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6742_2 ( .OUT(na6742_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6742_6 ( .RAM_O1(na6742_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6742_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x119y98     80'h00_0018_00_0000_0CEE_DA00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6743_1 ( .OUT(na6743_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na151_1), .IN6(1'b0), .IN7(~na102_1), .IN8(na92_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y70     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6744_4 ( .OUT(na6744_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2512_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6744_5 ( .OUT(na6744_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_109), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6744_6 ( .RAM_O2(na6744_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6744_2_i), .COMP_OUT(1'b0) );
// C_AND////      x113y63     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6745_1 ( .OUT(na6745_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na155_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y70     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6746_1 ( .OUT(na6746_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2510_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6746_2 ( .OUT(na6746_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_110), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6746_6 ( .RAM_O1(na6746_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6746_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y69     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6747_4 ( .OUT(na6747_2_i), .IN1(na2508_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6747_5 ( .OUT(na6747_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_111), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6747_6 ( .RAM_O2(na6747_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6747_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y69     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6748_1 ( .OUT(na6748_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2506_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6748_2 ( .OUT(na6748_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_112), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6748_6 ( .RAM_O1(na6748_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6748_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x99y100     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6749_1 ( .OUT(na6749_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na157_1), .IN7(~na2937_2), .IN8(na6750_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x86y90     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6750_1 ( .OUT(na6750_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9714_2), .IN5(~na1084_1), .IN6(1'b0), .IN7(~na920_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y68     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6751_4 ( .OUT(na6751_2_i), .IN1(na2504_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6751_5 ( .OUT(na6751_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_113), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6751_6 ( .RAM_O2(na6751_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6751_2_i), .COMP_OUT(1'b0) );
// C_OR////      x100y64     80'h00_0018_00_0000_0EEE_BE7D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6752_1 ( .OUT(na6752_1), .IN1(~na203_1), .IN2(na3718_1), .IN3(~na199_1), .IN4(~na6753_1), .IN5(na3720_2), .IN6(na3714_2),
                      .IN7(na9844_2), .IN8(~na207_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y60     80'h00_0018_00_0000_0888_4848
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6753_1 ( .OUT(na6753_1), .IN1(na186_1), .IN2(na182_1), .IN3(~na180_1), .IN4(na194_1), .IN5(na189_1), .IN6(na179_1), .IN7(~na180_2),
                      .IN8(na178_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y68     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6754_1 ( .OUT(na6754_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2502_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6754_2 ( .OUT(na6754_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_114), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6754_6 ( .RAM_O1(na6754_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6754_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y67     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6755_4 ( .OUT(na6755_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2500_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6755_5 ( .OUT(na6755_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_115), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6755_6 ( .RAM_O2(na6755_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6755_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y67     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6756_1 ( .OUT(na6756_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2498_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6756_2 ( .OUT(na6756_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_116), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6756_6 ( .RAM_O1(na6756_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6756_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y66     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6757_4 ( .OUT(na6757_2_i), .IN1(na2496_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6757_5 ( .OUT(na6757_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_117), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6757_6 ( .RAM_O2(na6757_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6757_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y66     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6758_1 ( .OUT(na6758_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2494_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6758_2 ( .OUT(na6758_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_118), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6758_6 ( .RAM_O1(na6758_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6758_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x81y78     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6759_1 ( .OUT(na6759_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na803_2), .IN6(~na2438_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y65     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6760_4 ( .OUT(na6760_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2492_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6760_5 ( .OUT(na6760_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_119), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6760_6 ( .RAM_O2(na6760_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6760_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y65     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6761_1 ( .OUT(na6761_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2490_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6761_2 ( .OUT(na6761_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6629_120), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6761_6 ( .RAM_O1(na6761_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6761_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x67y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6762_4 ( .OUT(na6762_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6762_6 ( .RAM_O2(na6762_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6762_2), .COMP_OUT(1'b0) );
// C_AND////      x67y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6763_1 ( .OUT(na6763_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6763_6 ( .RAM_O1(na6763_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6763_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x67y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6764_4 ( .OUT(na6764_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6764_6 ( .RAM_O2(na6764_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6764_2), .COMP_OUT(1'b0) );
// C_AND////      x67y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6765_1 ( .OUT(na6765_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6765_6 ( .RAM_O1(na6765_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6765_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x65y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6766_4 ( .OUT(na6766_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6766_6 ( .RAM_O2(na6766_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6766_2), .COMP_OUT(1'b0) );
// C_///XOR/      x87y75     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6767_4 ( .OUT(na6767_2), .IN1(1'b0), .IN2(na2962_1), .IN3(1'b0), .IN4(~na5585_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y78     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6768_1 ( .OUT(na6768_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1502_2), .IN8(~na2439_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y81     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6769_1 ( .OUT(na6769_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na9675_2), .IN5(~na2440_2), .IN6(1'b0), .IN7(~na807_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y77     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6770_1 ( .OUT(na6770_1), .IN1(1'b1), .IN2(na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na799_2), .IN6(~na2437_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x82y80     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6771_1 ( .OUT(na6771_1), .IN1(1'b1), .IN2(~na2773_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2443_2), .IN8(~na815_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6772_1 ( .OUT(na6772_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6772_6 ( .RAM_O1(na6772_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6772_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x65y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6773_4 ( .OUT(na6773_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6773_6 ( .RAM_O2(na6773_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6773_2), .COMP_OUT(1'b0) );
// C_MX2b////      x86y91     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6774_1 ( .OUT(na6774_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na9675_2), .IN5(~na811_2), .IN6(1'b0), .IN7(~na2441_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y80     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6775_1 ( .OUT(na6775_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na9675_2), .IN5(~na819_2), .IN6(1'b0), .IN7(~na2442_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x123y99     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6776_1 ( .OUT(na6776_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2951_2), .IN6(na6567_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x122y97     80'h00_0060_00_0000_0C0E_FF5A
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a6777_4 ( .OUT(na6777_2), .IN1(na8394_1), .IN2(1'b0), .IN3(~na755_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x123y98     80'h00_0078_00_0000_0C88_3C5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6778_1 ( .OUT(na6778_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6567_1), .IN7(1'b1), .IN8(~na2953_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6778_4 ( .OUT(na6778_2), .IN1(na6565_1), .IN2(1'b1), .IN3(~na709_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x126y98     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6779_4 ( .OUT(na6779_2), .IN1(~na6565_2), .IN2(1'b0), .IN3(1'b0), .IN4(na2953_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x128y99     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6780_4 ( .OUT(na6780_2), .IN1(1'b0), .IN2(na6563_1), .IN3(1'b0), .IN4(~na753_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x127y102     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6781_1 ( .OUT(na6781_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6565_1), .IN6(1'b1), .IN7(na709_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x127y102     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6782_4 ( .OUT(na6782_2), .IN1(1'b0), .IN2(na6563_2), .IN3(na709_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x125y101     80'h00_0018_00_0000_0CEE_A500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6783_1 ( .OUT(na6783_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na8394_1), .IN6(1'b0), .IN7(na755_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y101     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6784_1 ( .OUT(na6784_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na6567_1), .IN7(1'b1), .IN8(na2953_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6785_1 ( .OUT(na6785_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6785_6 ( .RAM_O1(na6785_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6785_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x94y104     80'h00_0018_00_0000_0888_8888
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6786_1 ( .OUT(na6786_1), .IN1(na251_1), .IN2(na252_1), .IN3(na3141_1), .IN4(na254_1), .IN5(na251_2), .IN6(na3148_1), .IN7(na3147_1),
                      .IN8(na3146_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y112     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6787_1 ( .OUT(na6787_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na291_2), .IN7(1'b1), .IN8(~na288_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y117     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6788_4 ( .OUT(na6788_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3906_1), .IN4(~na288_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y116     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6789_1 ( .OUT(na6789_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3906_2), .IN8(~na288_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y117     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6790_4 ( .OUT(na6790_2), .IN1(1'b1), .IN2(~na9191_2), .IN3(1'b1), .IN4(na3908_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y41     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6791_4 ( .OUT(na6791_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na2519_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6791_6 ( .RAM_O2(na6791_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6791_2), .COMP_OUT(1'b0) );
// C_///AND/      x129y67     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6792_4 ( .OUT(na6792_2), .IN1(~na296_1), .IN2(1'b1), .IN3(1'b1), .IN4(na295_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6793_4 ( .OUT(na6793_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6793_6 ( .RAM_O2(na6793_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6793_2), .COMP_OUT(1'b0) );
// C_OR////      x129y118     80'h00_0018_00_0000_0EEE_ACBC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6794_1 ( .OUT(na6794_1), .IN1(1'b0), .IN2(na318_1), .IN3(na320_2), .IN4(~na321_2), .IN5(1'b0), .IN6(na318_2), .IN7(na320_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6795_1 ( .OUT(na6795_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6795_6 ( .RAM_O1(na6795_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6795_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y115     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6796_4 ( .OUT(na6796_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na332_2), .IN4(~na9200_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y118     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6797_1 ( .OUT(na6797_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3899_1), .IN7(~na332_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y117     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6798_4 ( .OUT(na6798_2), .IN1(1'b1), .IN2(na3899_2), .IN3(~na332_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y117     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6799_1 ( .OUT(na6799_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3901_1), .IN6(1'b1), .IN7(~na332_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6800_4 ( .OUT(na6800_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6800_6 ( .RAM_O2(na6800_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6800_2), .COMP_OUT(1'b0) );
// C_AND////      x60y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6801_1 ( .OUT(na6801_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6801_6 ( .RAM_O1(na6801_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6801_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y46     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6802_4 ( .OUT(na6802_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2518_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6802_6 ( .RAM_O2(na6802_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6802_2), .COMP_OUT(1'b0) );
// C_AND////      x78y70     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6803_1 ( .OUT(na6803_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na356_1), .IN6(1'b1), .IN7(~na354_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y46     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6804_1 ( .OUT(na6804_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2517_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6804_6 ( .RAM_O1(na6804_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6804_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR////      x55y39     80'h00_0018_00_0000_0C66_C500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6805_1 ( .OUT(na6805_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2576_2), .IN6(1'b0), .IN7(1'b0), .IN8(na5685_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y45     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6806_4 ( .OUT(na6806_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2516_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6806_6 ( .RAM_O2(na6806_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6806_2), .COMP_OUT(1'b0) );
// C_///XOR/      x75y51     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6807_4 ( .OUT(na6807_2), .IN1(~na2574_2), .IN2(1'b0), .IN3(1'b0), .IN4(na5931_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y45     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6808_1 ( .OUT(na6808_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2515_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6808_6 ( .RAM_O1(na6808_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6808_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y44     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6809_4 ( .OUT(na6809_2), .IN1(na2514_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6809_6 ( .RAM_O2(na6809_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6809_2), .COMP_OUT(1'b0) );
// C_///AND/      x84y58     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6810_4 ( .OUT(na6810_2), .IN1(~na2566_1), .IN2(~na365_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6811_1 ( .OUT(na6811_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6811_6 ( .RAM_O1(na6811_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6811_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR////      x57y54     80'h00_0018_00_0000_0C66_C300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6812_1 ( .OUT(na6812_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na2586_2), .IN7(1'b0), .IN8(na5685_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y43     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6813_4 ( .OUT(na6813_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6813_6 ( .RAM_O2(na6813_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6813_2), .COMP_OUT(1'b0) );
// C_AND////      x60y43     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6814_1 ( .OUT(na6814_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6814_6 ( .RAM_O1(na6814_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6814_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6815_4 ( .OUT(na6815_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6815_6 ( .RAM_O2(na6815_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6815_2), .COMP_OUT(1'b0) );
// C_///OR/      x77y87     80'h00_0060_00_0000_0C0E_FFB3
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a6816_4 ( .OUT(na6816_2), .IN1(1'b0), .IN2(~na9246_2), .IN3(na3321_1), .IN4(~na3323_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6817_1 ( .OUT(na6817_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6817_6 ( .RAM_O1(na6817_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6817_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6818_4 ( .OUT(na6818_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6818_6 ( .RAM_O2(na6818_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6818_2), .COMP_OUT(1'b0) );
// C_AND////      x60y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6819_1 ( .OUT(na6819_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6819_6 ( .RAM_O1(na6819_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6819_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6820_4 ( .OUT(na6820_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6820_6 ( .RAM_O2(na6820_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6820_2), .COMP_OUT(1'b0) );
// C_AND////      x69y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6821_1 ( .OUT(na6821_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6821_6 ( .RAM_O1(na6821_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6821_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6822_4 ( .OUT(na6822_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6822_6 ( .RAM_O2(na6822_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6822_2), .COMP_OUT(1'b0) );
// C_MX4a////      x79y79     80'h00_0018_00_0040_0C86_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6823_1 ( .OUT(na6823_1), .IN1(1'b0), .IN2(na401_2), .IN3(na9211_2), .IN4(1'b1), .IN5(na402_1), .IN6(1'b1), .IN7(1'b1), .IN8(na341_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6824_1 ( .OUT(na6824_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6824_6 ( .RAM_O1(na6824_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6824_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y46     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6825_4 ( .OUT(na6825_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2582_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6825_6 ( .RAM_O2(na6825_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6825_2), .COMP_OUT(1'b0) );
// C_AND////      x69y46     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6826_1 ( .OUT(na6826_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2580_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6826_6 ( .RAM_O1(na6826_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6826_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y45     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6827_4 ( .OUT(na6827_2), .IN1(1'b1), .IN2(na2578_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6827_6 ( .RAM_O2(na6827_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6827_2), .COMP_OUT(1'b0) );
// C_AND////      x89y69     80'h00_0018_00_0000_0C88_15FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6828_1 ( .OUT(na6828_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na86_1), .IN6(1'b1), .IN7(~na66_1), .IN8(~na61_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y45     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6829_1 ( .OUT(na6829_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2576_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6829_6 ( .RAM_O1(na6829_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6829_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y44     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6830_4 ( .OUT(na6830_2), .IN1(na2574_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6830_6 ( .RAM_O2(na6830_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6830_2), .COMP_OUT(1'b0) );
// C_AND////      x69y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6831_1 ( .OUT(na6831_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6831_6 ( .RAM_O1(na6831_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6831_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y43     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6832_4 ( .OUT(na6832_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6832_6 ( .RAM_O2(na6832_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6832_2), .COMP_OUT(1'b0) );
// C_AND////      x69y43     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6833_1 ( .OUT(na6833_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6833_6 ( .RAM_O1(na6833_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6833_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x70y124     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6834_1 ( .OUT(na6834_1), .IN1(1'b1), .IN2(~na506_2), .IN3(1'b0), .IN4(1'b0), .IN5(na501_1), .IN6(na505_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6835_4 ( .OUT(na6835_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6835_6 ( .RAM_O2(na6835_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6835_2), .COMP_OUT(1'b0) );
// C_AND////      x71y89     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6836_1 ( .OUT(na6836_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na714_2), .IN6(na504_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6837_1 ( .OUT(na6837_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6837_6 ( .RAM_O1(na6837_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6837_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6838_4 ( .OUT(na6838_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6838_6 ( .RAM_O2(na6838_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6838_2), .COMP_OUT(1'b0) );
// C_AND///AND/      x77y88     80'h00_0078_00_0000_0C88_A8A2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6839_1 ( .OUT(na6839_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na514_2), .IN6(na504_1), .IN7(na517_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6839_4 ( .OUT(na6839_2), .IN1(na514_2), .IN2(~na504_1), .IN3(na517_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6840_1 ( .OUT(na6840_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6840_6 ( .RAM_O1(na6840_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6840_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x129y75     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6841_1 ( .OUT(na6841_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na515_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x62y48     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6842_4 ( .OUT(na6842_2_i), .IN1(na2488_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6842_5 ( .OUT(na6842_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6842_6 ( .RAM_O2(na6842_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6842_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y48     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6843_1 ( .OUT(na6843_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2486_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6843_2 ( .OUT(na6843_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6843_6 ( .RAM_O1(na6843_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6843_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y47     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6844_4 ( .OUT(na6844_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2484_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6844_5 ( .OUT(na6844_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6844_6 ( .RAM_O2(na6844_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6844_2_i), .COMP_OUT(1'b0) );
// C_///AND/      x68y85     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6845_4 ( .OUT(na6845_2), .IN1(na1373_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1407_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x62y47     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6846_1 ( .OUT(na6846_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2480_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6846_2 ( .OUT(na6846_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6846_6 ( .RAM_O1(na6846_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6846_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x77y85     80'h00_0018_00_0000_0EEE_0BD3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6847_1 ( .OUT(na6847_1), .IN1(1'b0), .IN2(~na3325_1), .IN3(~na517_1), .IN4(na406_1), .IN5(na353_1), .IN6(~na396_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y48     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6848_4 ( .OUT(na6848_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2477_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6848_5 ( .OUT(na6848_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6848_6 ( .RAM_O2(na6848_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6848_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x67y120     80'h00_0018_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6849_1 ( .OUT(na6849_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na531_2), .IN8(~na527_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y48     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6850_1 ( .OUT(na6850_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2474_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6850_2 ( .OUT(na6850_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6850_6 ( .RAM_O1(na6850_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6850_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y47     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6851_4 ( .OUT(na6851_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2471_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6851_5 ( .OUT(na6851_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6851_6 ( .RAM_O2(na6851_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6851_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y47     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6852_1 ( .OUT(na6852_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2468_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6852_2 ( .OUT(na6852_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6852_6 ( .RAM_O1(na6852_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6852_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///ORAND/      x72y84     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a6853_4 ( .OUT(na6853_2), .IN1(~na3305_1), .IN2(~na9439_2), .IN3(~na3308_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y46     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6854_4 ( .OUT(na6854_2_i), .IN1(1'b1), .IN2(na2465_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6854_5 ( .OUT(na6854_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6854_6 ( .RAM_O2(na6854_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6854_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x70y118     80'h00_0018_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6855_1 ( .OUT(na6855_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na531_1), .IN8(~na532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y46     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6856_1 ( .OUT(na6856_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2462_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6856_2 ( .OUT(na6856_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6856_6 ( .RAM_O1(na6856_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6856_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y45     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6857_4 ( .OUT(na6857_2_i), .IN1(1'b1), .IN2(na2459_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6857_5 ( .OUT(na6857_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6857_6 ( .RAM_O2(na6857_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6857_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y45     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6858_1 ( .OUT(na6858_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2455_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6858_2 ( .OUT(na6858_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6858_6 ( .RAM_O1(na6858_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6858_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x78y82     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6859_1 ( .OUT(na6859_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3305_1), .IN6(~na3107_2), .IN7(~na3308_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y44     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6860_4 ( .OUT(na6860_2_i), .IN1(1'b1), .IN2(na2454_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6860_5 ( .OUT(na6860_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6860_6 ( .RAM_O2(na6860_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6860_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y44     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6861_1 ( .OUT(na6861_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3583_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6861_2 ( .OUT(na6861_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6861_6 ( .RAM_O1(na6861_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6861_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y43     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6862_4 ( .OUT(na6862_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3580_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6862_5 ( .OUT(na6862_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6862_6 ( .RAM_O2(na6862_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6862_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y43     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6863_1 ( .OUT(na6863_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3577_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6863_2 ( .OUT(na6863_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6863_6 ( .RAM_O1(na6863_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6863_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x78y79     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6864_1 ( .OUT(na6864_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3305_1), .IN6(~na9348_2), .IN7(~na3308_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y42     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6865_4 ( .OUT(na6865_2_i), .IN1(1'b1), .IN2(na3574_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6865_5 ( .OUT(na6865_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6865_6 ( .RAM_O2(na6865_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6865_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x66y120     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6866_1 ( .OUT(na6866_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na546_2), .IN6(na536_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x66y87     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6867_1 ( .OUT(na6867_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2177_1), .IN6(~na9818_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x74y86     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6868_4 ( .OUT(na6868_2), .IN1(1'b1), .IN2(na5459_1), .IN3(1'b1), .IN4(na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x71y116     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a6869_4 ( .OUT(na6869_2), .IN1(~na2256_1), .IN2(~na9817_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x71y111     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6870_1 ( .OUT(na6870_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1373_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3319_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y122     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6871_1 ( .OUT(na6871_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na542_1), .IN8(na9257_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y42     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6872_1 ( .OUT(na6872_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3571_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6872_2 ( .OUT(na6872_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6872_6 ( .RAM_O1(na6872_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6872_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y41     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6873_4 ( .OUT(na6873_2_i), .IN1(na3568_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6873_5 ( .OUT(na6873_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6873_6 ( .RAM_O2(na6873_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6873_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y41     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6874_1 ( .OUT(na6874_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3565_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6874_2 ( .OUT(na6874_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6874_6 ( .RAM_O1(na6874_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6874_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x63y117     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6875_1 ( .OUT(na6875_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9260_2), .IN8(na551_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y46     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6876_4 ( .OUT(na6876_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2512_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6876_5 ( .OUT(na6876_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_89), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6876_6 ( .RAM_O2(na6876_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6876_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y46     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6877_1 ( .OUT(na6877_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2510_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6877_2 ( .OUT(na6877_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_90), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6877_6 ( .RAM_O1(na6877_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6877_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y45     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6878_4 ( .OUT(na6878_2_i), .IN1(na2508_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6878_5 ( .OUT(na6878_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_91), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6878_6 ( .RAM_O2(na6878_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6878_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x57y122     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6879_1 ( .OUT(na6879_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9263_2), .IN8(na557_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y45     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6880_1 ( .OUT(na6880_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2506_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6880_2 ( .OUT(na6880_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_92), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6880_6 ( .RAM_O1(na6880_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6880_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x103y95     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6881_4 ( .OUT(na6881_2), .IN1(na1860_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na896_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y44     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6882_4 ( .OUT(na6882_2_i), .IN1(na2504_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6882_5 ( .OUT(na6882_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_93), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6882_6 ( .RAM_O2(na6882_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6882_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y44     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6883_1 ( .OUT(na6883_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2502_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6883_2 ( .OUT(na6883_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_94), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6883_6 ( .RAM_O1(na6883_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6883_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y43     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6884_4 ( .OUT(na6884_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2500_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6884_5 ( .OUT(na6884_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_95), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6884_6 ( .RAM_O2(na6884_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6884_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y43     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6885_1 ( .OUT(na6885_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2498_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6885_2 ( .OUT(na6885_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_96), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6885_6 ( .RAM_O1(na6885_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6885_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x59y122     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6886_1 ( .OUT(na6886_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9269_2), .IN8(na578_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x72y97     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6887_1 ( .OUT(na6887_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1379_2), .IN8(na3309_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x65y112     80'h00_0078_00_0000_0CEE_3370
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a6888_1 ( .OUT(na6888_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3317_1), .IN7(1'b0), .IN8(~na587_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a6888_4 ( .OUT(na6888_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na3308_1), .IN4(~na587_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x66y108     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6889_4 ( .OUT(na6889_2), .IN1(1'b1), .IN2(1'b1), .IN3(na5463_1), .IN4(na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y42     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6890_4 ( .OUT(na6890_2_i), .IN1(na2496_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6890_5 ( .OUT(na6890_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_97), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6890_6 ( .RAM_O2(na6890_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6890_2_i), .COMP_OUT(1'b0) );
// C_///AND/      x55y125     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6891_4 ( .OUT(na6891_2), .IN1(na2185_1), .IN2(na9818_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x58y124     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6892_1 ( .OUT(na6892_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na9271_2), .IN6(na582_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y42     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6893_1 ( .OUT(na6893_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2494_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6893_2 ( .OUT(na6893_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_98), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6893_6 ( .RAM_O1(na6893_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6893_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y41     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6894_4 ( .OUT(na6894_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2492_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6894_5 ( .OUT(na6894_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_99), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6894_6 ( .RAM_O2(na6894_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6894_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y41     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6895_1 ( .OUT(na6895_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2490_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a6895_2 ( .OUT(na6895_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6630_100), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6895_6 ( .RAM_O1(na6895_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6895_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x52y124     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6896_1 ( .OUT(na6896_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9273_2), .IN8(na592_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6897_4 ( .OUT(na6897_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6897_6 ( .RAM_O2(na6897_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6897_2), .COMP_OUT(1'b0) );
// C_AND////      x67y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6898_1 ( .OUT(na6898_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6898_6 ( .RAM_O1(na6898_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6898_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x67y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6899_4 ( .OUT(na6899_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6899_6 ( .RAM_O2(na6899_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6899_2), .COMP_OUT(1'b0) );
// C_MX2b////      x52y122     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6900_1 ( .OUT(na6900_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9277_2), .IN8(na593_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6901_1 ( .OUT(na6901_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6901_6 ( .RAM_O1(na6901_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6901_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x65y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6902_4 ( .OUT(na6902_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6902_6 ( .RAM_O2(na6902_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6902_2), .COMP_OUT(1'b0) );
// C_AND////      x65y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6903_1 ( .OUT(na6903_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6903_6 ( .RAM_O1(na6903_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6903_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x58y123     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6904_1 ( .OUT(na6904_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9279_2), .IN8(na602_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6905_4 ( .OUT(na6905_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6905_6 ( .RAM_O2(na6905_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6905_2), .COMP_OUT(1'b0) );
// C_AND////      x65y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6906_1 ( .OUT(na6906_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6906_6 ( .RAM_O1(na6906_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6906_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x99y1     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6907_1 ( .OUT(na6907_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6907_6 ( .RAM_O1(na6907_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6907_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y8     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6908_4 ( .OUT(na6908_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6908_6 ( .RAM_O2(na6908_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6908_2), .COMP_OUT(1'b0) );
// C_MX2b////      x53y124     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6909_1 ( .OUT(na6909_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na608_1), .IN8(na603_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y8     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6910_1 ( .OUT(na6910_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6910_6 ( .RAM_O1(na6910_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6910_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y7     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6911_4 ( .OUT(na6911_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6911_6 ( .RAM_O2(na6911_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6911_2), .COMP_OUT(1'b0) );
// C_AND////      x92y7     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6912_1 ( .OUT(na6912_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6912_6 ( .RAM_O1(na6912_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6912_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x53y121     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6913_1 ( .OUT(na6913_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9283_2), .IN8(na613_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y6     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6914_4 ( .OUT(na6914_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6914_6 ( .RAM_O2(na6914_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6914_2), .COMP_OUT(1'b0) );
// C_AND////      x92y6     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6915_1 ( .OUT(na6915_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6915_6 ( .RAM_O1(na6915_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6915_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y5     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6916_4 ( .OUT(na6916_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6916_6 ( .RAM_O2(na6916_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6916_2), .COMP_OUT(1'b0) );
// C_MX2b////      x57y119     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6917_1 ( .OUT(na6917_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9285_2), .IN8(na618_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y5     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6918_1 ( .OUT(na6918_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6918_6 ( .RAM_O1(na6918_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6918_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y4     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6919_4 ( .OUT(na6919_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6919_6 ( .RAM_O2(na6919_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6919_2), .COMP_OUT(1'b0) );
// C_AND////      x92y4     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6920_1 ( .OUT(na6920_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6920_6 ( .RAM_O1(na6920_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6920_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x59y123     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6921_1 ( .OUT(na6921_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9288_2), .IN8(na623_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y3     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6922_4 ( .OUT(na6922_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6922_6 ( .RAM_O2(na6922_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6922_2), .COMP_OUT(1'b0) );
// C_AND////      x92y3     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6923_1 ( .OUT(na6923_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6923_6 ( .RAM_O1(na6923_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6923_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y2     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6924_4 ( .OUT(na6924_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6924_6 ( .RAM_O2(na6924_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6924_2), .COMP_OUT(1'b0) );
// C_MX2b////      x61y118     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6925_1 ( .OUT(na6925_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9291_2), .IN8(na628_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y2     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6926_1 ( .OUT(na6926_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6926_6 ( .RAM_O1(na6926_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6926_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y1     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6927_4 ( .OUT(na6927_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6927_6 ( .RAM_O2(na6927_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6927_2), .COMP_OUT(1'b0) );
// C_AND////      x92y1     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6928_1 ( .OUT(na6928_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6928_6 ( .RAM_O1(na6928_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6928_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x59y121     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6929_1 ( .OUT(na6929_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9293_2), .IN8(na629_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y3     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6930_4 ( .OUT(na6930_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6930_6 ( .RAM_O2(na6930_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6930_2), .COMP_OUT(1'b0) );
// C_AND////      x101y3     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6931_1 ( .OUT(na6931_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6931_6 ( .RAM_O1(na6931_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6931_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y2     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6932_4 ( .OUT(na6932_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6932_6 ( .RAM_O2(na6932_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6932_2), .COMP_OUT(1'b0) );
// C_MX2b////      x51y124     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6933_1 ( .OUT(na6933_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9295_2), .IN8(na638_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y2     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6934_1 ( .OUT(na6934_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6934_6 ( .RAM_O1(na6934_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6934_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x121y95     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6935_1 ( .OUT(na6935_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na643_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2953_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x135y93     80'h00_0078_00_0000_0C88_53A4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6936_1 ( .OUT(na6936_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2894_2), .IN7(~na3546_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6936_4 ( .OUT(na6936_2), .IN1(~na7054_2), .IN2(na2919_1), .IN3(na106_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x135y74     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6937_4 ( .OUT(na6937_2), .IN1(~na3542_1), .IN2(1'b1), .IN3(~na2838_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x127y95     80'h00_0018_00_0040_0A16_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6938_1 ( .OUT(na6938_1), .IN1(1'b1), .IN2(na2894_2), .IN3(1'b1), .IN4(na2836_2), .IN5(na7054_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y1     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6939_4 ( .OUT(na6939_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6939_6 ( .RAM_O2(na6939_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6939_2), .COMP_OUT(1'b0) );
// C_AND////      x101y1     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6940_1 ( .OUT(na6940_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6940_6 ( .RAM_O1(na6940_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6940_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x96y3     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6941_2 ( .OUT(na6941_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6631_36), .CP_O(1'b0) );
// C_MX2b////      x67y118     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6942_1 ( .OUT(na6942_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9300_2), .IN8(na662_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x96y2     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6943_5 ( .OUT(na6943_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6631_37), .CP_O(1'b0) );
// C_/RAM_I1///      x96y2     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6944_2 ( .OUT(na6944_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6631_38), .CP_O(1'b0) );
// C_////RAM_I2      x96y1     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6945_5 ( .OUT(na6945_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6631_39), .CP_O(1'b0) );
// C_MX2b////      x65y119     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6946_1 ( .OUT(na6946_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9304_2), .IN8(na668_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x96y1     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6947_2 ( .OUT(na6947_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6631_40), .CP_O(1'b0) );
// C_AND////      x131y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6948_1 ( .OUT(na6948_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6948_6 ( .RAM_O1(na6948_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6948_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y88     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6949_4 ( .OUT(na6949_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6949_6 ( .RAM_O2(na6949_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6949_2), .COMP_OUT(1'b0) );
// C_MX2b////      x57y123     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6950_1 ( .OUT(na6950_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9305_2), .IN8(na669_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y88     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6951_1 ( .OUT(na6951_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6951_6 ( .RAM_O1(na6951_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6951_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y87     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6952_4 ( .OUT(na6952_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6952_6 ( .RAM_O2(na6952_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6952_2), .COMP_OUT(1'b0) );
// C_AND////      x124y87     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6953_1 ( .OUT(na6953_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6953_6 ( .RAM_O1(na6953_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6953_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x61y119     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6954_1 ( .OUT(na6954_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9306_2), .IN8(na674_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y86     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6955_4 ( .OUT(na6955_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6955_6 ( .RAM_O2(na6955_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6955_2), .COMP_OUT(1'b0) );
// C_AND////      x124y86     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6956_1 ( .OUT(na6956_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6956_6 ( .RAM_O1(na6956_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6956_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y85     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6957_4 ( .OUT(na6957_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6957_6 ( .RAM_O2(na6957_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6957_2), .COMP_OUT(1'b0) );
// C_MX2b////      x59y124     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6958_1 ( .OUT(na6958_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9308_2), .IN8(na683_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y85     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6959_1 ( .OUT(na6959_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6959_6 ( .RAM_O1(na6959_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6959_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y84     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6960_4 ( .OUT(na6960_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6960_6 ( .RAM_O2(na6960_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6960_2), .COMP_OUT(1'b0) );
// C_AND////      x124y84     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6961_1 ( .OUT(na6961_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6961_6 ( .RAM_O1(na6961_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6961_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x64y122     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6962_1 ( .OUT(na6962_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9309_2), .IN8(na688_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y83     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6963_4 ( .OUT(na6963_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6963_6 ( .RAM_O2(na6963_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6963_2), .COMP_OUT(1'b0) );
// C_AND////      x124y83     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6964_1 ( .OUT(na6964_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6964_6 ( .RAM_O1(na6964_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6964_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y82     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6965_4 ( .OUT(na6965_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6965_6 ( .RAM_O2(na6965_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6965_2), .COMP_OUT(1'b0) );
// C_MX2b////      x55y123     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6966_1 ( .OUT(na6966_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9312_2), .IN8(na693_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6967_1 ( .OUT(na6967_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6967_6 ( .RAM_O1(na6967_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6967_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6968_4 ( .OUT(na6968_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6968_6 ( .RAM_O2(na6968_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6968_2), .COMP_OUT(1'b0) );
// C_AND////      x124y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6969_1 ( .OUT(na6969_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6969_6 ( .RAM_O1(na6969_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6969_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x63y120     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6970_1 ( .OUT(na6970_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9314_2), .IN8(na698_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x133y83     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6971_4 ( .OUT(na6971_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6971_6 ( .RAM_O2(na6971_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6971_2), .COMP_OUT(1'b0) );
// C_AND////      x133y83     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6972_1 ( .OUT(na6972_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6972_6 ( .RAM_O1(na6972_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6972_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y82     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6973_4 ( .OUT(na6973_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6973_6 ( .RAM_O2(na6973_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6973_2), .COMP_OUT(1'b0) );
// C_MX2b////      x61y120     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6974_1 ( .OUT(na6974_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9317_2), .IN8(na703_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6975_1 ( .OUT(na6975_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6975_6 ( .RAM_O1(na6975_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6975_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6976_4 ( .OUT(na6976_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6976_6 ( .RAM_O2(na6976_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6976_2), .COMP_OUT(1'b0) );
// C_AND////      x133y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6977_1 ( .OUT(na6977_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6977_6 ( .RAM_O1(na6977_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6977_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x65y120     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6978_1 ( .OUT(na6978_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9319_2), .IN8(na704_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x128y83     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6979_2 ( .OUT(na6979_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6632_36), .CP_O(1'b0) );
// C_AND////      x121y94     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6980_1 ( .OUT(na6980_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na643_1), .IN6(1'b1), .IN7(na709_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x128y82     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6981_5 ( .OUT(na6981_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6632_37), .CP_O(1'b0) );
// C_/RAM_I1///      x128y82     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6982_2 ( .OUT(na6982_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6632_38), .CP_O(1'b0) );
// C_////RAM_I2      x128y81     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6983_5 ( .OUT(na6983_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6632_39), .CP_O(1'b0) );
// C_/RAM_I1///      x128y81     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a6984_2 ( .OUT(na6984_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6632_40), .CP_O(1'b0) );
// C_AND////      x99y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6985_1 ( .OUT(na6985_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6985_6 ( .RAM_O1(na6985_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6985_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y104     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6986_4 ( .OUT(na6986_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6986_6 ( .RAM_O2(na6986_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6986_2), .COMP_OUT(1'b0) );
// C_AND////      x92y104     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6987_1 ( .OUT(na6987_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6987_6 ( .RAM_O1(na6987_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6987_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x57y124     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6988_1 ( .OUT(na6988_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9322_2), .IN8(na724_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y103     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6989_4 ( .OUT(na6989_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6989_6 ( .RAM_O2(na6989_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6989_2), .COMP_OUT(1'b0) );
// C_AND////      x67y91     80'h00_0018_00_0000_0C88_C4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6990_1 ( .OUT(na6990_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na714_1), .IN6(na727_2), .IN7(1'b1), .IN8(na725_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y103     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6991_1 ( .OUT(na6991_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6991_6 ( .RAM_O1(na6991_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6991_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x77y93     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6992_1 ( .OUT(na6992_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na740_2), .IN6(na728_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y102     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6993_4 ( .OUT(na6993_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6993_6 ( .RAM_O2(na6993_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na6993_2), .COMP_OUT(1'b0) );
// C_AND////      x92y102     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6994_1 ( .OUT(na6994_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a6994_6 ( .RAM_O1(na6994_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na6994_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x121y98     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6995_4 ( .OUT(na6995_2), .IN1(na643_1), .IN2(1'b1), .IN3(na709_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y100     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6996_1 ( .OUT(na6996_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na740_1), .IN6(na737_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x62y98     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6997_1 ( .OUT(na6997_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na741_1), .IN6(na748_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y88     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6998_1 ( .OUT(na6998_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na745_1), .IN6(na748_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y99     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a6999_1 ( .OUT(na6999_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na749_1), .IN6(na1555_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y101     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7000_4 ( .OUT(na7000_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7000_6 ( .RAM_O2(na7000_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7000_2), .COMP_OUT(1'b0) );
// C_AND////      x123y95     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7001_1 ( .OUT(na7001_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na643_1), .IN6(1'b1), .IN7(1'b1), .IN8(na753_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y101     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7002_1 ( .OUT(na7002_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7002_6 ( .RAM_O1(na7002_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7002_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x121y98     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7003_1 ( .OUT(na7003_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na643_1), .IN6(1'b1), .IN7(na755_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x89y89     80'h00_0060_00_0000_0C0E_FFB5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7004_4 ( .OUT(na7004_2), .IN1(~na2960_1), .IN2(1'b0), .IN3(na757_1), .IN4(~na783_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y100     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7005_4 ( .OUT(na7005_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7005_6 ( .RAM_O2(na7005_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7005_2), .COMP_OUT(1'b0) );
// C_MX2b////      x65y100     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7006_1 ( .OUT(na7006_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na766_2), .IN6(na759_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y100     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7007_1 ( .OUT(na7007_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na766_1), .IN6(na763_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y98     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7008_1 ( .OUT(na7008_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na774_2), .IN8(na767_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y98     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7009_1 ( .OUT(na7009_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na774_1), .IN8(na771_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x69y115     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7010_1 ( .OUT(na7010_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na782_2), .IN8(na775_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x61y94     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7011_1 ( .OUT(na7011_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na782_1), .IN8(na779_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y100     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7012_1 ( .OUT(na7012_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7012_6 ( .RAM_O1(na7012_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7012_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y99     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7013_4 ( .OUT(na7013_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7013_6 ( .RAM_O2(na7013_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7013_2), .COMP_OUT(1'b0) );
// C_MX2b////      x66y100     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7014_1 ( .OUT(na7014_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na795_2), .IN6(na786_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y115     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7015_1 ( .OUT(na7015_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na795_1), .IN6(na792_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y99     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7016_1 ( .OUT(na7016_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7016_6 ( .RAM_O1(na7016_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7016_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x79y94     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7017_1 ( .OUT(na7017_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9338_2), .IN8(na806_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y99     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7018_1 ( .OUT(na7018_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9339_2), .IN8(na806_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y95     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7019_1 ( .OUT(na7019_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na807_1), .IN8(na810_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y102     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7020_1 ( .OUT(na7020_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na811_1), .IN6(na822_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y99     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7021_1 ( .OUT(na7021_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na826_2), .IN8(na815_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y97     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7022_1 ( .OUT(na7022_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na819_1), .IN6(na822_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y100     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7023_1 ( .OUT(na7023_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na826_1), .IN8(na823_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y100     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7024_1 ( .OUT(na7024_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na828_1), .IN8(na831_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x78y100     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7025_1 ( .OUT(na7025_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1497_2), .IN8(na834_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y101     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7026_1 ( .OUT(na7026_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na860_2), .IN6(na843_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y101     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7027_1 ( .OUT(na7027_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na866_2), .IN8(na847_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x107y96     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7028_1 ( .OUT(na7028_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2253_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y95     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7029_1 ( .OUT(na7029_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3118_1), .IN6(na9345_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y98     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7030_4 ( .OUT(na7030_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7030_6 ( .RAM_O2(na7030_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7030_2), .COMP_OUT(1'b0) );
// C_MX2b////      x66y101     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7031_1 ( .OUT(na7031_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na860_1), .IN6(na857_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x107y103     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7032_1 ( .OUT(na7032_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na8_2), .IN8(~na2761_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x103y92     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7033_4 ( .OUT(na7033_2), .IN1(na853_2), .IN2(1'b1), .IN3(na3113_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y102     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7034_1 ( .OUT(na7034_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na866_1), .IN8(na863_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y98     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7035_1 ( .OUT(na7035_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7035_6 ( .RAM_O1(na7035_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7035_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x117y69     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7036_1 ( .OUT(na7036_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na981_1), .IN7(1'b1), .IN8(~na839_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y97     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7037_4 ( .OUT(na7037_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7037_6 ( .RAM_O2(na7037_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7037_2), .COMP_OUT(1'b0) );
// C_///OR/      x115y105     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7038_4 ( .OUT(na7038_2), .IN1(~na481_1), .IN2(1'b0), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y110     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7039_1 ( .OUT(na7039_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3119_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x107y94     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7040_4 ( .OUT(na7040_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na8_2), .IN4(~na2716_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y107     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7041_1 ( .OUT(na7041_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(na3170_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x101y92     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7042_4 ( .OUT(na7042_2), .IN1(~na9133_2), .IN2(1'b0), .IN3(~na1116_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y95     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7043_4 ( .OUT(na7043_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3192_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x123y70     80'h00_0060_00_0000_0C0E_FF75
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7044_4 ( .OUT(na7044_2), .IN1(~na900_1), .IN2(1'b0), .IN3(~na1119_1), .IN4(~na1333_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7045_1 ( .OUT(na7045_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7045_6 ( .RAM_O1(na7045_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7045_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x105y97     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7046_1 ( .OUT(na7046_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3161_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y110     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7047_1 ( .OUT(na7047_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2721_1), .IN6(na9345_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y99     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7048_4 ( .OUT(na7048_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7048_6 ( .RAM_O2(na7048_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7048_2), .COMP_OUT(1'b0) );
// C_///AND/      x75y100     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7049_4 ( .OUT(na7049_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na4853_2), .IN4(na2155_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y99     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7050_1 ( .OUT(na7050_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7050_6 ( .RAM_O1(na7050_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7050_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR////      x119y97     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7051_1 ( .OUT(na7051_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1064_1), .IN7(na9369_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x130y45     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7052_4 ( .OUT(na7052_2), .IN1(~na9372_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y98     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7053_4 ( .OUT(na7053_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7053_6 ( .RAM_O2(na7053_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7053_2), .COMP_OUT(1'b0) );
// C_AND///AND/      x125y99     80'h00_0078_00_0000_0C88_1F52
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7054_1 ( .OUT(na7054_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2838_1), .IN8(~na2836_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7054_4 ( .OUT(na7054_2), .IN1(na995_1), .IN2(~na2671_1), .IN3(~na2673_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x126y97     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7055_1 ( .OUT(na7055_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2838_1), .IN8(na2836_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y98     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7056_1 ( .OUT(na7056_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7056_6 ( .RAM_O1(na7056_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7056_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///XOR/      x111y93     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7057_4 ( .OUT(na7057_2), .IN1(na1006_2), .IN2(na1007_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y97     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7058_4 ( .OUT(na7058_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7058_6 ( .RAM_O2(na7058_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7058_2), .COMP_OUT(1'b0) );
// C_XOR////      x130y61     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7059_1 ( .OUT(na7059_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1008_2), .IN7(1'b0), .IN8(na1009_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7060_1 ( .OUT(na7060_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7060_6 ( .RAM_O1(na7060_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7060_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x96y99     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7061_2 ( .OUT(na7061_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6633_36), .CP_O(1'b0) );
// C_///XOR/      x118y78     80'h00_0060_00_0000_0C06_FFAA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7062_4 ( .OUT(na7062_2), .IN1(na1020_1), .IN2(1'b0), .IN3(na1021_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y104     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7063_1 ( .OUT(na7063_1), .IN1(~na853_2), .IN2(~na9486_2), .IN3(~na8_2), .IN4(~na4897_2), .IN5(~na9487_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x96y98     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7064_5 ( .OUT(na7064_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6633_37), .CP_O(1'b0) );
// C_/RAM_I1///      x96y98     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7065_2 ( .OUT(na7065_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6633_38), .CP_O(1'b0) );
// C_////RAM_I2      x96y97     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7066_5 ( .OUT(na7066_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6633_39), .CP_O(1'b0) );
// C_/RAM_I1///      x96y97     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7067_2 ( .OUT(na7067_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6633_40), .CP_O(1'b0) );
// C_AND////      x79y61     80'h00_0018_00_0000_0C88_23FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7068_1 ( .OUT(na7068_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na35_1), .IN7(na432_1), .IN8(~na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7069_1 ( .OUT(na7069_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7069_6 ( .RAM_O1(na7069_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7069_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y88     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7070_4 ( .OUT(na7070_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7070_6 ( .RAM_O2(na7070_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7070_2), .COMP_OUT(1'b0) );
// C_AND////      x129y76     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7071_1 ( .OUT(na7071_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1048_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x93y99     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7072_1 ( .OUT(na7072_1), .IN1(~na853_2), .IN2(~na9653_2), .IN3(~na8_2), .IN4(~na4900_2), .IN5(~na9654_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y88     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7073_1 ( .OUT(na7073_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7073_6 ( .RAM_O1(na7073_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7073_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y87     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7074_4 ( .OUT(na7074_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7074_6 ( .RAM_O2(na7074_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7074_2), .COMP_OUT(1'b0) );
// C_AND////      x92y87     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7075_1 ( .OUT(na7075_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7075_6 ( .RAM_O1(na7075_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7075_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x118y75     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7076_1 ( .OUT(na7076_1), .IN1(~na488_1), .IN2(~na3011_1), .IN3(~na8_2), .IN4(~na2168_1), .IN5(~na3114_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y86     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7077_4 ( .OUT(na7077_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7077_6 ( .RAM_O2(na7077_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7077_2), .COMP_OUT(1'b0) );
// C_OR////      x107y69     80'h00_0018_00_0000_0EEE_CEBA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7078_1 ( .OUT(na7078_1), .IN1(na488_1), .IN2(1'b0), .IN3(na567_1), .IN4(~na856_2), .IN5(na1028_1), .IN6(na955_1), .IN7(1'b0),
                      .IN8(na9352_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y86     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7079_1 ( .OUT(na7079_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7079_6 ( .RAM_O1(na7079_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7079_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y85     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7080_4 ( .OUT(na7080_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7080_6 ( .RAM_O2(na7080_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7080_2), .COMP_OUT(1'b0) );
// C_AND////      x92y85     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7081_1 ( .OUT(na7081_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7081_6 ( .RAM_O1(na7081_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7081_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x120y83     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7082_1 ( .OUT(na7082_1), .IN1(~na488_1), .IN2(~na3010_1), .IN3(~na8_2), .IN4(~na2968_1), .IN5(~na3121_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y84     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7083_4 ( .OUT(na7083_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7083_6 ( .RAM_O2(na7083_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7083_2), .COMP_OUT(1'b0) );
// C_AND////      x92y84     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7084_1 ( .OUT(na7084_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7084_6 ( .RAM_O1(na7084_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7084_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y83     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7085_4 ( .OUT(na7085_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7085_6 ( .RAM_O2(na7085_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7085_2), .COMP_OUT(1'b0) );
// C_ORAND////      x120y75     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7086_1 ( .OUT(na7086_1), .IN1(~na488_1), .IN2(~na3009_1), .IN3(~na8_2), .IN4(~na3066_1), .IN5(~na1658_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y83     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7087_1 ( .OUT(na7087_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7087_6 ( .RAM_O1(na7087_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7087_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y82     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7088_4 ( .OUT(na7088_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7088_6 ( .RAM_O2(na7088_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7088_2), .COMP_OUT(1'b0) );
// C_AND////      x92y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7089_1 ( .OUT(na7089_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7089_6 ( .RAM_O1(na7089_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7089_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x130y46     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7090_1 ( .OUT(na7090_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3888_1), .IN8(~na989_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7091_4 ( .OUT(na7091_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7091_6 ( .RAM_O2(na7091_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7091_2), .COMP_OUT(1'b0) );
// C_AND////      x92y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7092_1 ( .OUT(na7092_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7092_6 ( .RAM_O1(na7092_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7092_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y83     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7093_4 ( .OUT(na7093_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7093_6 ( .RAM_O2(na7093_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7093_2), .COMP_OUT(1'b0) );
// C_AND////      x129y74     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7094_1 ( .OUT(na7094_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1128_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y83     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7095_1 ( .OUT(na7095_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7095_6 ( .RAM_O1(na7095_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7095_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x109y58     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7096_1 ( .OUT(na7096_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9413_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y58     80'h00_0018_00_0000_0CEE_0D00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7097_1 ( .OUT(na7097_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2991_1), .IN6(na974_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y57     80'h00_0018_00_0000_0888_1F15
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7098_1 ( .OUT(na7098_1), .IN1(~na1167_1), .IN2(1'b1), .IN3(~na1165_2), .IN4(~na1134_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na1165_1),
                      .IN8(~na1134_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y82     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7099_4 ( .OUT(na7099_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7099_6 ( .RAM_O2(na7099_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7099_2), .COMP_OUT(1'b0) );
// C_AND////      x125y71     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7100_1 ( .OUT(na7100_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7101_1 ( .OUT(na7101_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7101_6 ( .RAM_O1(na7101_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7101_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x127y63     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7102_4 ( .OUT(na7102_2), .IN1(~na296_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1142_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7103_4 ( .OUT(na7103_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7103_6 ( .RAM_O2(na7103_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7103_2), .COMP_OUT(1'b0) );
// C_AND////      x101y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7104_1 ( .OUT(na7104_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7104_6 ( .RAM_O1(na7104_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7104_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x96y83     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7105_2 ( .OUT(na7105_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6634_36), .CP_O(1'b0) );
// C_AND////      x109y56     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7106_1 ( .OUT(na7106_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1167_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x96y82     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7107_5 ( .OUT(na7107_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6634_37), .CP_O(1'b0) );
// C_AND////      x85y94     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7108_1 ( .OUT(na7108_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1177_2), .IN8(na9440_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y86     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7109_1 ( .OUT(na7109_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1224_1), .IN6(na1173_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x96y82     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7110_2 ( .OUT(na7110_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6634_38), .CP_O(1'b0) );
// C_AND////      x87y95     80'h00_0018_00_0000_0888_1555
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7111_1 ( .OUT(na7111_1), .IN1(~na1193_1), .IN2(1'b1), .IN3(~na1191_2), .IN4(1'b1), .IN5(~na1193_2), .IN6(1'b1), .IN7(~na1191_1),
                      .IN8(~na1188_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x96y81     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7112_5 ( .OUT(na7112_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6634_39), .CP_O(1'b0) );
// C_/RAM_I1///      x96y81     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7113_2 ( .OUT(na7113_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6634_40), .CP_O(1'b0) );
// C_///AND/      x85y93     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7114_4 ( .OUT(na7114_2), .IN1(1'b1), .IN2(na1189_2), .IN3(1'b1), .IN4(na1188_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7115_1 ( .OUT(na7115_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7115_6 ( .RAM_O1(na7115_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7115_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y40     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7116_4 ( .OUT(na7116_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7116_6 ( .RAM_O2(na7116_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7116_2), .COMP_OUT(1'b0) );
// C_AND////      x28y40     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7117_1 ( .OUT(na7117_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7117_6 ( .RAM_O1(na7117_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7117_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x87y96     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7118_1 ( .OUT(na7118_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1193_1), .IN6(na1189_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y39     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7119_4 ( .OUT(na7119_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7119_6 ( .RAM_O2(na7119_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7119_2), .COMP_OUT(1'b0) );
// C_///AND/      x87y91     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7120_4 ( .OUT(na7120_2), .IN1(na1193_2), .IN2(na1189_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y39     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7121_1 ( .OUT(na7121_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7121_6 ( .RAM_O1(na7121_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7121_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x89y93     80'h00_0078_00_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7122_1 ( .OUT(na7122_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1189_2), .IN7(na1191_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7122_4 ( .OUT(na7122_2), .IN1(1'b1), .IN2(na1189_2), .IN3(na1191_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y38     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7123_4 ( .OUT(na7123_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7123_6 ( .RAM_O2(na7123_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7123_2), .COMP_OUT(1'b0) );
// C_AND////      x99y112     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7124_1 ( .OUT(na7124_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1900_1), .IN6(1'b1), .IN7(na1275_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y38     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7125_1 ( .OUT(na7125_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7125_6 ( .RAM_O1(na7125_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7125_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7126_4 ( .OUT(na7126_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7126_6 ( .RAM_O2(na7126_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7126_2), .COMP_OUT(1'b0) );
// C_AND////      x28y37     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7127_1 ( .OUT(na7127_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7127_6 ( .RAM_O1(na7127_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7127_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y36     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7128_4 ( .OUT(na7128_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7128_6 ( .RAM_O2(na7128_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7128_2), .COMP_OUT(1'b0) );
// C_MX2b////      x51y122     80'h00_0018_00_0040_0AA8_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7129_1 ( .OUT(na7129_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1380_1), .IN5(1'b0), .IN6(na582_1), .IN7(1'b0), .IN8(~na1381_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y36     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7130_1 ( .OUT(na7130_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7130_6 ( .RAM_O1(na7130_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7130_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x77y50     80'h00_0018_00_0000_0888_5531
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7131_1 ( .OUT(na7131_1), .IN1(~na2562_1), .IN2(~na2561_1), .IN3(1'b1), .IN4(~na2563_1), .IN5(~na2559_1), .IN6(1'b1), .IN7(~na2560_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y60     80'h00_0060_00_0000_0C08_FFA1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7132_4 ( .OUT(na7132_2), .IN1(~na2565_1), .IN2(~na2564_1), .IN3(na2558_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y112     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7133_1 ( .OUT(na7133_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na503_2), .IN5(1'b0), .IN6(na3977_1), .IN7(1'b0), .IN8(na3980_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x62y120     80'h00_0018_00_0040_0A51_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7134_1 ( .OUT(na7134_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1380_1), .IN5(~na1389_1), .IN6(1'b0), .IN7(na542_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x55y121     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7135_1 ( .OUT(na7135_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1388_1), .IN6(1'b1), .IN7(na359_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x120y85     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7136_1 ( .OUT(na7136_1), .IN1(~na488_1), .IN2(~na2915_1), .IN3(~na8_2), .IN4(~na1382_1), .IN5(~na3196_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y35     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7137_4 ( .OUT(na7137_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7137_6 ( .RAM_O2(na7137_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7137_2), .COMP_OUT(1'b0) );
// C_AND////      x28y35     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7138_1 ( .OUT(na7138_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7138_6 ( .RAM_O1(na7138_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7138_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y34     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7139_4 ( .OUT(na7139_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7139_6 ( .RAM_O2(na7139_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7139_2), .COMP_OUT(1'b0) );
// C_MX2b////      x76y114     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7140_1 ( .OUT(na7140_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na503_2), .IN5(na3979_1), .IN6(1'b0), .IN7(na3982_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x67y111     80'h00_0078_00_0000_0CEE_3533
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7141_1 ( .OUT(na7141_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1403_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na3309_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7141_4 ( .OUT(na7141_2), .IN1(1'b0), .IN2(~na3317_1), .IN3(1'b0), .IN4(~na1399_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y110     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7142_4 ( .OUT(na7142_2), .IN1(1'b1), .IN2(na5467_2), .IN3(1'b1), .IN4(na3309_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7143_1 ( .OUT(na7143_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7143_6 ( .RAM_O1(na7143_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7143_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x72y83     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7144_4 ( .OUT(na7144_2), .IN1(1'b1), .IN2(na3259_1), .IN3(1'b1), .IN4(na3319_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x67y116     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7145_1 ( .OUT(na7145_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1620_1), .IN6(1'b0), .IN7(~na3308_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x62y116     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7146_4 ( .OUT(na7146_2), .IN1(na3313_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2193_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y116     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7147_1 ( .OUT(na7147_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1400_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1393_1), .IN7(1'b0), .IN8(na1399_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x118y87     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7148_1 ( .OUT(na7148_1), .IN1(~na488_1), .IN2(~na2914_1), .IN3(~na8_2), .IN4(~na832_1), .IN5(~na3203_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7149_4 ( .OUT(na7149_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7149_6 ( .RAM_O2(na7149_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7149_2), .COMP_OUT(1'b0) );
// C_AND////      x28y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7150_1 ( .OUT(na7150_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7150_6 ( .RAM_O1(na7150_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7150_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7151_4 ( .OUT(na7151_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7151_6 ( .RAM_O2(na7151_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7151_2), .COMP_OUT(1'b0) );
// C_AND////      x59y116     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7152_1 ( .OUT(na7152_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9280_2), .IN6(na1393_1), .IN7(1'b1), .IN8(na1380_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7153_1 ( .OUT(na7153_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7153_6 ( .RAM_O1(na7153_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7153_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x56y119     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7154_1 ( .OUT(na7154_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1403_1), .IN6(1'b1), .IN7(na359_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7155_4 ( .OUT(na7155_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7155_6 ( .RAM_O2(na7155_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7155_2), .COMP_OUT(1'b0) );
// C_AND////      x37y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7156_1 ( .OUT(na7156_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7156_6 ( .RAM_O1(na7156_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7156_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x74y85     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7157_4 ( .OUT(na7157_2), .IN1(~na1405_1), .IN2(1'b1), .IN3(na359_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y117     80'h00_0018_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7158_1 ( .OUT(na7158_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1400_1), .IN4(1'b1), .IN5(na9503_2), .IN6(1'b0), .IN7(na542_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7159_4 ( .OUT(na7159_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7159_6 ( .RAM_O2(na7159_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7159_2), .COMP_OUT(1'b0) );
// C_MX2b////      x114y57     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7160_1 ( .OUT(na7160_1), .IN1(1'b1), .IN2(na9463_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1409_1), .IN8(~na6447_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x111y86     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7161_1 ( .OUT(na7161_1), .IN1(~na488_1), .IN2(~na3110_1), .IN3(~na8_2), .IN4(~na3070_1), .IN5(~na2239_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7162_1 ( .OUT(na7162_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7162_6 ( .RAM_O1(na7162_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7162_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_////RAM_I2      x32y34     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7163_5 ( .OUT(na7163_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6635_37), .CP_O(1'b0) );
// C_/RAM_I1///      x32y34     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7164_2 ( .OUT(na7164_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6635_38), .CP_O(1'b0) );
// C_ORAND////      x110y99     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7165_1 ( .OUT(na7165_1), .IN1(~na488_1), .IN2(~na1270_1), .IN3(~na8_2), .IN4(~na1207_1), .IN5(~na1104_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x32y33     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7166_5 ( .OUT(na7166_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6635_39), .CP_O(1'b0) );
// C_/RAM_I1///      x32y33     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7167_2 ( .OUT(na7167_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6635_40), .CP_O(1'b0) );
// C_AND////      x35y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7168_1 ( .OUT(na7168_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7168_6 ( .RAM_O1(na7168_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7168_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y104     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7169_4 ( .OUT(na7169_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7169_6 ( .RAM_O2(na7169_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7169_2), .COMP_OUT(1'b0) );
// C_AND////      x28y104     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7170_1 ( .OUT(na7170_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7170_6 ( .RAM_O1(na7170_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7170_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x108y84     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7171_1 ( .OUT(na7171_1), .IN1(~na853_2), .IN2(~na2780_1), .IN3(~na567_1), .IN4(~na2710_1), .IN5(~na9684_2), .IN6(~na1042_1),
                      .IN7(~na1033_1), .IN8(~na9242_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y103     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7172_4 ( .OUT(na7172_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7172_6 ( .RAM_O2(na7172_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7172_2), .COMP_OUT(1'b0) );
// C_AND////      x28y103     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7173_1 ( .OUT(na7173_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7173_6 ( .RAM_O1(na7173_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7173_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y102     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7174_4 ( .OUT(na7174_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7174_6 ( .RAM_O2(na7174_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7174_2), .COMP_OUT(1'b0) );
// C_AND////      x28y102     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7175_1 ( .OUT(na7175_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7175_6 ( .RAM_O1(na7175_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7175_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x118y43     80'h00_0018_00_0000_0EEE_C5EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7176_1 ( .OUT(na7176_1), .IN1(na1427_1), .IN2(1'b0), .IN3(na9508_2), .IN4(na1429_2), .IN5(~na1430_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na1429_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y101     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7177_4 ( .OUT(na7177_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7177_6 ( .RAM_O2(na7177_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7177_2), .COMP_OUT(1'b0) );
// C_ORAND////      x118y80     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7178_1 ( .OUT(na7178_1), .IN1(~na488_1), .IN2(~na486_1), .IN3(~na567_1), .IN4(~na2708_1), .IN5(~na2793_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y101     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7179_1 ( .OUT(na7179_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7179_6 ( .RAM_O1(na7179_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7179_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y100     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7180_4 ( .OUT(na7180_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7180_6 ( .RAM_O2(na7180_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7180_2), .COMP_OUT(1'b0) );
// C_AND////      x28y100     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7181_1 ( .OUT(na7181_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7181_6 ( .RAM_O1(na7181_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7181_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x110y96     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7182_4 ( .OUT(na7182_2), .IN1(~na941_1), .IN2(~na1042_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y101     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7183_1 ( .OUT(na7183_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6012_1), .IN6(1'b1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x120y98     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7184_4 ( .OUT(na7184_2), .IN1(1'b0), .IN2(~na1042_1), .IN3(1'b0), .IN4(~na940_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y105     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7185_1 ( .OUT(na7185_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9133_2), .IN6(1'b1), .IN7(na6011_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x108y94     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7186_4 ( .OUT(na7186_2), .IN1(1'b0), .IN2(~na1042_1), .IN3(1'b0), .IN4(~na939_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x114y105     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7187_1 ( .OUT(na7187_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6010_1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x106y94     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7188_4 ( .OUT(na7188_2), .IN1(~na938_1), .IN2(~na1042_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y105     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7189_1 ( .OUT(na7189_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9133_2), .IN6(1'b1), .IN7(na6009_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x114y91     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7190_1 ( .OUT(na7190_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na937_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x116y102     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7191_1 ( .OUT(na7191_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9133_2), .IN6(1'b1), .IN7(na6008_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x116y99     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7192_1 ( .OUT(na7192_1), .IN1(~na2693_1), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na6007_2), .IN5(~na936_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y99     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7193_4 ( .OUT(na7193_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7193_6 ( .RAM_O2(na7193_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7193_2), .COMP_OUT(1'b0) );
// C_AND////      x28y99     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7194_1 ( .OUT(na7194_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7194_6 ( .RAM_O1(na7194_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7194_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y98     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7195_4 ( .OUT(na7195_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7195_6 ( .RAM_O2(na7195_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7195_2), .COMP_OUT(1'b0) );
// C_AND////      x28y98     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7196_1 ( .OUT(na7196_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7196_6 ( .RAM_O1(na7196_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7196_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y97     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7197_4 ( .OUT(na7197_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7197_6 ( .RAM_O2(na7197_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7197_2), .COMP_OUT(1'b0) );
// C_ORAND////      x116y100     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7198_1 ( .OUT(na7198_1), .IN1(~na1870_1), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na6006_1), .IN5(~na935_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7199_1 ( .OUT(na7199_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7199_6 ( .RAM_O1(na7199_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7199_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y99     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7200_4 ( .OUT(na7200_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7200_6 ( .RAM_O2(na7200_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7200_2), .COMP_OUT(1'b0) );
// C_AND////      x37y99     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7201_1 ( .OUT(na7201_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7201_6 ( .RAM_O1(na7201_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7201_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x125y103     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7202_4 ( .OUT(na7202_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2734_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x115y108     80'h00_0078_00_0000_0CEE_7053
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7203_1 ( .OUT(na7203_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na8_2), .IN8(~na6005_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7203_4 ( .OUT(na7203_2), .IN1(1'b0), .IN2(~na1042_1), .IN3(~na933_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y105     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7204_1 ( .OUT(na7204_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na488_1), .IN6(1'b1), .IN7(na930_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y98     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7205_4 ( .OUT(na7205_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7205_6 ( .RAM_O2(na7205_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7205_2), .COMP_OUT(1'b0) );
// C_///AND/      x126y75     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7206_4 ( .OUT(na7206_2), .IN1(na1039_1), .IN2(na955_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x60y119     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7207_1 ( .OUT(na7207_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1400_1), .IN4(1'b1), .IN5(1'b0), .IN6(na582_1), .IN7(1'b0), .IN8(na587_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y92     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7208_1 ( .OUT(na7208_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na428_1), .IN6(1'b1), .IN7(~na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x100y80     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7209_1 ( .OUT(na7209_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(~na2699_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y81     80'h00_0078_00_0000_0C88_ACA4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7210_1 ( .OUT(na7210_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6590_1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7210_4 ( .OUT(na7210_2), .IN1(~na9166_2), .IN2(na89_1), .IN3(na8_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y111     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7211_1 ( .OUT(na7211_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na503_2), .IN5(1'b0), .IN6(na3977_2), .IN7(1'b0), .IN8(na3980_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7212_1 ( .OUT(na7212_1), .IN1(~na488_1), .IN2(~na9490_2), .IN3(~na567_1), .IN4(~na1128_2), .IN5(~na2790_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y98     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7213_1 ( .OUT(na7213_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7213_6 ( .RAM_O1(na7213_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7213_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y97     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7214_4 ( .OUT(na7214_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7214_6 ( .RAM_O2(na7214_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7214_2), .COMP_OUT(1'b0) );
// C_AND////      x37y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7215_1 ( .OUT(na7215_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7215_6 ( .RAM_O1(na7215_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7215_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x115y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7216_1 ( .OUT(na7216_1), .IN1(~na488_1), .IN2(~na9396_2), .IN3(~na567_1), .IN4(~na295_1), .IN5(~na9683_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x32y99     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7217_2 ( .OUT(na7217_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6636_36), .CP_O(1'b0) );
// C_////RAM_I2      x32y98     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7218_5 ( .OUT(na7218_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6636_37), .CP_O(1'b0) );
// C_/RAM_I1///      x32y98     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7219_2 ( .OUT(na7219_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6636_38), .CP_O(1'b0) );
// C_ORAND////      x122y80     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7220_1 ( .OUT(na7220_1), .IN1(~na488_1), .IN2(~na2701_1), .IN3(~na567_1), .IN4(~na515_1), .IN5(~na2741_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x32y97     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7221_5 ( .OUT(na7221_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6636_39), .CP_O(1'b0) );
// C_/RAM_I1///      x32y97     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7222_2 ( .OUT(na7222_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6636_40), .CP_O(1'b0) );
// C_AND////      x131y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7223_1 ( .OUT(na7223_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7223_6 ( .RAM_O1(na7223_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7223_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x118y86     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7224_1 ( .OUT(na7224_1), .IN1(~na488_1), .IN2(~na892_1), .IN3(~na567_1), .IN4(~na1048_2), .IN5(~na2792_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y72     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7225_4 ( .OUT(na7225_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7225_6 ( .RAM_O2(na7225_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7225_2), .COMP_OUT(1'b0) );
// C_AND////      x124y72     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7226_1 ( .OUT(na7226_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7226_6 ( .RAM_O1(na7226_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7226_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y71     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7227_4 ( .OUT(na7227_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7227_6 ( .RAM_O2(na7227_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7227_2), .COMP_OUT(1'b0) );
// C_ORAND////      x117y106     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7228_1 ( .OUT(na7228_1), .IN1(~na488_1), .IN2(~na9662_2), .IN3(~na567_1), .IN4(~na2706_2), .IN5(~na2794_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y71     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7229_1 ( .OUT(na7229_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7229_6 ( .RAM_O1(na7229_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7229_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y70     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7230_4 ( .OUT(na7230_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7230_6 ( .RAM_O2(na7230_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7230_2), .COMP_OUT(1'b0) );
// C_AND////      x124y70     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7231_1 ( .OUT(na7231_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7231_6 ( .RAM_O1(na7231_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7231_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x71y103     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7232_1 ( .OUT(na7232_1), .IN1(na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1497_1), .IN8(na1494_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y102     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7233_1 ( .OUT(na7233_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1498_1), .IN8(na831_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y93     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7234_1 ( .OUT(na7234_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1502_1), .IN8(na810_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x110y88     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7235_1 ( .OUT(na7235_1), .IN1(~na853_2), .IN2(~na9669_2), .IN3(~na567_1), .IN4(~na2712_1), .IN5(~na2796_1), .IN6(~na1042_1),
                      .IN7(~na9241_2), .IN8(~na9663_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y69     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7236_4 ( .OUT(na7236_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7236_6 ( .RAM_O2(na7236_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7236_2), .COMP_OUT(1'b0) );
// C_AND////      x124y69     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7237_1 ( .OUT(na7237_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7237_6 ( .RAM_O1(na7237_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7237_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y68     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7238_4 ( .OUT(na7238_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7238_6 ( .RAM_O2(na7238_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7238_2), .COMP_OUT(1'b0) );
// C_AND////      x124y68     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7239_1 ( .OUT(na7239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7239_6 ( .RAM_O1(na7239_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7239_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x115y83     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7240_1 ( .OUT(na7240_1), .IN1(~na853_2), .IN2(~na2781_1), .IN3(~na567_1), .IN4(~na1142_1), .IN5(~na2743_1), .IN6(~na1042_1),
                      .IN7(~na2704_1), .IN8(~na9242_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y67     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7241_4 ( .OUT(na7241_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7241_6 ( .RAM_O2(na7241_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7241_2), .COMP_OUT(1'b0) );
// C_AND////      x124y67     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7242_1 ( .OUT(na7242_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7242_6 ( .RAM_O1(na7242_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7242_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y66     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7243_4 ( .OUT(na7243_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7243_6 ( .RAM_O2(na7243_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7243_2), .COMP_OUT(1'b0) );
// C_AND////      x124y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7244_1 ( .OUT(na7244_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7244_6 ( .RAM_O1(na7244_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7244_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x110y80     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7245_1 ( .OUT(na7245_1), .IN1(~na853_2), .IN2(~na2782_1), .IN3(~na567_1), .IN4(~na1140_1), .IN5(~na9670_2), .IN6(~na1042_1),
                      .IN7(~na1123_1), .IN8(~na9242_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7246_4 ( .OUT(na7246_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7246_6 ( .RAM_O2(na7246_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7246_2), .COMP_OUT(1'b0) );
// C_AND////      x124y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7247_1 ( .OUT(na7247_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7247_6 ( .RAM_O1(na7247_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7247_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y67     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7248_4 ( .OUT(na7248_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7248_6 ( .RAM_O2(na7248_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7248_2), .COMP_OUT(1'b0) );
// C_AND////      x133y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7249_1 ( .OUT(na7249_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7249_6 ( .RAM_O1(na7249_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7249_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x108y80     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7250_1 ( .OUT(na7250_1), .IN1(~na853_2), .IN2(~na2783_1), .IN3(~na567_1), .IN4(~na2714_1), .IN5(~na9685_2), .IN6(~na1042_1),
                      .IN7(~na9241_2), .IN8(~na1121_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x133y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7251_4 ( .OUT(na7251_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7251_6 ( .RAM_O2(na7251_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7251_2), .COMP_OUT(1'b0) );
// C_AND////      x133y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7252_1 ( .OUT(na7252_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7252_6 ( .RAM_O1(na7252_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7252_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7253_4 ( .OUT(na7253_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7253_6 ( .RAM_O2(na7253_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7253_2), .COMP_OUT(1'b0) );
// C_AND////      x133y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7254_1 ( .OUT(na7254_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7254_6 ( .RAM_O1(na7254_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7254_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x109y80     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7255_1 ( .OUT(na7255_1), .IN1(~na853_2), .IN2(~na2784_1), .IN3(~na567_1), .IN4(~na2774_1), .IN5(~na2764_1), .IN6(~na1042_1),
                      .IN7(~na1118_1), .IN8(~na9242_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x128y67     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7256_2 ( .OUT(na7256_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6637_36), .CP_O(1'b0) );
// C_////RAM_I2      x128y66     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7257_5 ( .OUT(na7257_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6637_37), .CP_O(1'b0) );
// C_/RAM_I1///      x128y66     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7258_2 ( .OUT(na7258_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6637_38), .CP_O(1'b0) );
// C_////RAM_I2      x128y65     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7259_5 ( .OUT(na7259_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6637_39), .CP_O(1'b0) );
// C_OR////      x97y78     80'h00_0018_00_0000_0EEE_E30B
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7260_1 ( .OUT(na7260_1), .IN1(na7265_1), .IN2(~na7262_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na7262_1), .IN7(na7263_2),
                      .IN8(na1531_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x128y65     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7261_2 ( .OUT(na7261_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6637_40), .CP_O(1'b0) );
// C_OR///OR/      x97y80     80'h00_0078_00_0000_0CEE_3333
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7262_1 ( .OUT(na7262_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1524_1), .IN7(1'b0), .IN8(~na2776_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7262_4 ( .OUT(na7262_2), .IN1(1'b0), .IN2(~na1042_1), .IN3(1'b0), .IN4(~na2801_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y79     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7263_4 ( .OUT(na7263_2), .IN1(na9519_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2785_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x131y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7264_1 ( .OUT(na7264_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7264_6 ( .RAM_O1(na7264_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7264_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x101y87     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7265_1 ( .OUT(na7265_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1530_1), .IN8(na1117_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x113y80     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7266_1 ( .OUT(na7266_1), .IN1(~na853_2), .IN2(~na2786_1), .IN3(~na567_1), .IN4(~na2778_1), .IN5(~na2802_1), .IN6(~na1042_1),
                      .IN7(~na9241_2), .IN8(~na2705_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y56     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7267_4 ( .OUT(na7267_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7267_6 ( .RAM_O2(na7267_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7267_2), .COMP_OUT(1'b0) );
// C_AND////      x124y56     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7268_1 ( .OUT(na7268_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7268_6 ( .RAM_O1(na7268_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7268_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y55     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7269_4 ( .OUT(na7269_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7269_6 ( .RAM_O2(na7269_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7269_2), .COMP_OUT(1'b0) );
// C_AND////      x124y55     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7270_1 ( .OUT(na7270_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7270_6 ( .RAM_O1(na7270_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7270_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x112y78     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7271_1 ( .OUT(na7271_1), .IN1(~na853_2), .IN2(~na9682_2), .IN3(~na567_1), .IN4(~na2723_2), .IN5(~na2803_1), .IN6(~na1042_1),
                      .IN7(~na9405_2), .IN8(~na9242_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y54     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7272_4 ( .OUT(na7272_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7272_6 ( .RAM_O2(na7272_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7272_2), .COMP_OUT(1'b0) );
// C_AND////      x124y54     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7273_1 ( .OUT(na7273_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7273_6 ( .RAM_O1(na7273_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7273_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y53     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7274_4 ( .OUT(na7274_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7274_6 ( .RAM_O2(na7274_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7274_2), .COMP_OUT(1'b0) );
// C_AND////      x124y53     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7275_1 ( .OUT(na7275_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7275_6 ( .RAM_O1(na7275_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7275_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x116y78     80'h00_0018_00_0000_0888_54F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7276_1 ( .OUT(na7276_1), .IN1(~na7277_2), .IN2(na7278_2), .IN3(1'b1), .IN4(1'b1), .IN5(~na7279_1), .IN6(na7278_1), .IN7(~na7281_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x121y73     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7277_4 ( .OUT(na7277_2), .IN1(1'b1), .IN2(na99_2), .IN3(1'b1), .IN4(na9362_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x109y88     80'h00_0078_00_0000_0CEE_5355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7278_1 ( .OUT(na7278_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(~na2804_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7278_4 ( .OUT(na7278_2), .IN1(~na488_1), .IN2(1'b0), .IN3(~na1114_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x115y73     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7279_1 ( .OUT(na7279_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9266_2), .IN6(1'b1), .IN7(na2735_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y52     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7280_4 ( .OUT(na7280_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7280_6 ( .RAM_O2(na7280_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7280_2), .COMP_OUT(1'b0) );
// C_///AND/      x110y91     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7281_4 ( .OUT(na7281_2), .IN1(na853_2), .IN2(1'b1), .IN3(na2787_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x123y97     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7282_1 ( .OUT(na7282_1), .IN1(~na853_2), .IN2(~na9689_2), .IN3(~na8_2), .IN4(~na4919_2), .IN5(~na9690_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y52     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7283_1 ( .OUT(na7283_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7283_6 ( .RAM_O1(na7283_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7283_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y51     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7284_4 ( .OUT(na7284_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7284_6 ( .RAM_O2(na7284_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7284_2), .COMP_OUT(1'b0) );
// C_AND////      x124y51     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7285_1 ( .OUT(na7285_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7285_6 ( .RAM_O1(na7285_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7285_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x108y87     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7286_1 ( .OUT(na7286_1), .IN1(~na853_2), .IN2(~na9687_2), .IN3(~na8_2), .IN4(~na4917_2), .IN5(~na9688_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y50     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7287_4 ( .OUT(na7287_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7287_6 ( .RAM_O2(na7287_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7287_2), .COMP_OUT(1'b0) );
// C_AND////      x124y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7288_1 ( .OUT(na7288_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7288_6 ( .RAM_O1(na7288_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7288_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7289_4 ( .OUT(na7289_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7289_6 ( .RAM_O2(na7289_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7289_2), .COMP_OUT(1'b0) );
// C_OR////      x116y73     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7290_1 ( .OUT(na7290_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na882_1), .IN6(~na1042_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x126y76     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7291_4 ( .OUT(na7291_2), .IN1(na869_1), .IN2(1'b1), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x112y72     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7292_1 ( .OUT(na7292_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na881_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y71     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7293_1 ( .OUT(na7293_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na868_1), .IN6(1'b1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y114     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7294_1 ( .OUT(na7294_1), .IN1(~na734_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1552_1), .IN6(na1555_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x118y72     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7295_4 ( .OUT(na7295_2), .IN1(1'b0), .IN2(~na1042_1), .IN3(1'b0), .IN4(~na880_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x122y71     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7296_1 ( .OUT(na7296_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na867_1), .IN6(1'b1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x116y67     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7297_4 ( .OUT(na7297_2), .IN1(~na879_1), .IN2(~na1042_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x128y74     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7298_4 ( .OUT(na7298_2), .IN1(na480_1), .IN2(1'b1), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x118y71     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7299_4 ( .OUT(na7299_2), .IN1(1'b0), .IN2(~na1042_1), .IN3(1'b0), .IN4(~na1893_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x118y72     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7300_1 ( .OUT(na7300_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na479_1), .IN6(1'b1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y68     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7301_1 ( .OUT(na7301_1), .IN1(~na1127_1), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na883_1), .IN5(~na9539_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7302_1 ( .OUT(na7302_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7302_6 ( .RAM_O1(na7302_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7302_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y51     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7303_4 ( .OUT(na7303_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7303_6 ( .RAM_O2(na7303_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7303_2), .COMP_OUT(1'b0) );
// C_AND////      x133y51     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7304_1 ( .OUT(na7304_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7304_6 ( .RAM_O1(na7304_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7304_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x123y73     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7305_1 ( .OUT(na7305_1), .IN1(~na9370_2), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na1367_1), .IN5(~na877_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x133y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7306_4 ( .OUT(na7306_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7306_6 ( .RAM_O2(na7306_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7306_2), .COMP_OUT(1'b0) );
// C_AND////      x133y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7307_1 ( .OUT(na7307_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7307_6 ( .RAM_O1(na7307_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7307_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7308_4 ( .OUT(na7308_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7308_6 ( .RAM_O2(na7308_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7308_2), .COMP_OUT(1'b0) );
// C_AND////      x133y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7309_1 ( .OUT(na7309_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7309_6 ( .RAM_O1(na7309_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7309_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x114y74     80'h00_0018_00_0000_0888_CC51
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7310_1 ( .OUT(na7310_1), .IN1(~na3594_1), .IN2(~na3356_1), .IN3(~na3219_1), .IN4(1'b1), .IN5(1'b1), .IN6(na3555_1), .IN7(1'b1),
                      .IN8(na9362_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x108y65     80'h00_0078_00_0000_0CEE_5570
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7311_1 ( .OUT(na7311_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na853_2), .IN6(1'b0), .IN7(~na1895_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7311_4 ( .OUT(na7311_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na567_1), .IN4(~na870_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y68     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7312_4 ( .OUT(na7312_2), .IN1(na906_1), .IN2(1'b1), .IN3(na904_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7313_1 ( .OUT(na7313_1), .IN1(~na853_2), .IN2(~na9691_2), .IN3(~na8_2), .IN4(~na4922_2), .IN5(~na9692_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x128y51     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7314_2 ( .OUT(na7314_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6638_36), .CP_O(1'b0) );
// C_////RAM_I2      x128y50     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7315_5 ( .OUT(na7315_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6638_37), .CP_O(1'b0) );
// C_/RAM_I1///      x128y50     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7316_2 ( .OUT(na7316_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6638_38), .CP_O(1'b0) );
// C_OR////      x100y95     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7317_1 ( .OUT(na7317_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na895_1), .IN6(~na1042_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x102y104     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7318_4 ( .OUT(na7318_2), .IN1(1'b1), .IN2(na560_1), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x112y86     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7319_1 ( .OUT(na7319_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na1366_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y105     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7320_4 ( .OUT(na7320_2), .IN1(1'b1), .IN2(na1898_1), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x104y97     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7321_1 ( .OUT(na7321_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na1364_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y98     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7322_1 ( .OUT(na7322_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1363_1), .IN6(1'b1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x98y87     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7323_1 ( .OUT(na7323_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na902_1), .IN6(~na1042_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x106y102     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7324_4 ( .OUT(na7324_2), .IN1(na1362_1), .IN2(1'b1), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x102y91     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7325_1 ( .OUT(na7325_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na897_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y102     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7326_1 ( .OUT(na7326_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1899_1), .IN6(1'b1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x110y106     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7327_1 ( .OUT(na7327_1), .IN1(~na313_1), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na9494_2), .IN5(~na9350_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x128y49     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7328_5 ( .OUT(na7328_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6638_39), .CP_O(1'b0) );
// C_/RAM_I1///      x128y49     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7329_2 ( .OUT(na7329_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6638_40), .CP_O(1'b0) );
// C_AND////      x131y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7330_1 ( .OUT(na7330_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7330_6 ( .RAM_O1(na7330_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7330_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y40     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7331_4 ( .OUT(na7331_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7331_6 ( .RAM_O2(na7331_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7331_2), .COMP_OUT(1'b0) );
// C_AND////      x124y40     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7332_1 ( .OUT(na7332_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7332_6 ( .RAM_O1(na7332_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7332_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y39     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7333_4 ( .OUT(na7333_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7333_6 ( .RAM_O2(na7333_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7333_2), .COMP_OUT(1'b0) );
// C_MX2b////      x63y118     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7334_1 ( .OUT(na7334_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9521_2), .IN8(na1587_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x122y93     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7335_1 ( .OUT(na7335_1), .IN1(~na1860_1), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na1353_1), .IN5(~na1897_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y39     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7336_1 ( .OUT(na7336_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7336_6 ( .RAM_O1(na7336_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7336_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y38     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7337_4 ( .OUT(na7337_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7337_6 ( .RAM_O2(na7337_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7337_2), .COMP_OUT(1'b0) );
// C_AND////      x124y38     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7338_1 ( .OUT(na7338_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7338_6 ( .RAM_O1(na7338_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7338_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x85y97     80'h00_0018_00_0000_0EEE_7EDA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7339_1 ( .OUT(na7339_1), .IN1(na7345_1), .IN2(1'b0), .IN3(~na7344_1), .IN4(na7343_2), .IN5(na7345_2), .IN6(na7347_1), .IN7(~na7344_2),
                      .IN8(~na7346_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7340_4 ( .OUT(na7340_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7340_6 ( .RAM_O2(na7340_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7340_2), .COMP_OUT(1'b0) );
// C_AND////      x124y37     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7341_1 ( .OUT(na7341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7341_6 ( .RAM_O1(na7341_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7341_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y36     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7342_4 ( .OUT(na7342_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7342_6 ( .RAM_O2(na7342_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7342_2), .COMP_OUT(1'b0) );
// C_///AND/      x100y98     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7343_4 ( .OUT(na7343_2), .IN1(na1860_1), .IN2(1'b1), .IN3(na9241_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x90y101     80'h00_0078_00_0000_0CEE_3555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7344_1 ( .OUT(na7344_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na906_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1346_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7344_4 ( .OUT(na7344_2), .IN1(~na428_1), .IN2(1'b0), .IN3(~na568_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x85y95     80'h00_0078_00_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7345_1 ( .OUT(na7345_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1524_1), .IN7(na561_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7345_4 ( .OUT(na7345_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1344_2), .IN4(na1527_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x86y96     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7346_1 ( .OUT(na7346_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1350_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1531_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x93y90     80'h00_0018_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7347_1 ( .OUT(na7347_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na285_1), .IN6(~na7348_1), .IN7(na9523_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x91y92     80'h00_0018_00_0000_0EEE_EDAC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7348_1 ( .OUT(na7348_1), .IN1(1'b0), .IN2(na3299_2), .IN3(na3276_1), .IN4(1'b0), .IN5(~na3588_1), .IN6(na3424_2), .IN7(na3301_1),
                      .IN8(na3216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y36     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7349_1 ( .OUT(na7349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7349_6 ( .RAM_O1(na7349_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7349_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y35     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7350_4 ( .OUT(na7350_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7350_6 ( .RAM_O2(na7350_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7350_2), .COMP_OUT(1'b0) );
// C_AND////      x124y35     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7351_1 ( .OUT(na7351_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7351_6 ( .RAM_O1(na7351_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7351_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y34     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7352_4 ( .OUT(na7352_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7352_6 ( .RAM_O2(na7352_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7352_2), .COMP_OUT(1'b0) );
// C_MX2b////      x58y121     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7353_1 ( .OUT(na7353_1), .IN1(~na526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9525_2), .IN8(na1604_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x96y88     80'h00_0018_00_0000_0888_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7354_1 ( .OUT(na7354_1), .IN1(~na488_1), .IN2(~na9438_2), .IN3(~na1177_1), .IN4(~na9362_2), .IN5(~na10164_2), .IN6(~na1042_1),
                      .IN7(~na567_1), .IN8(~na9476_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7355_1 ( .OUT(na7355_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7355_6 ( .RAM_O1(na7355_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7355_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7356_4 ( .OUT(na7356_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7356_6 ( .RAM_O2(na7356_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7356_2), .COMP_OUT(1'b0) );
// C_AND////      x124y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7357_1 ( .OUT(na7357_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7357_6 ( .RAM_O1(na7357_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7357_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7358_4 ( .OUT(na7358_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7358_6 ( .RAM_O2(na7358_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7358_2), .COMP_OUT(1'b0) );
// C_OR///OR/      x90y67     80'h00_0078_00_0000_0CEE_B00B
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7359_1 ( .OUT(na7359_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1177_1), .IN8(~na1527_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7359_4 ( .OUT(na7359_2), .IN1(na2991_1), .IN2(~na1612_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y89     80'h00_0018_00_0000_0888_5544
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7360_1 ( .OUT(na7360_1), .IN1(~na1193_2), .IN2(na1614_1), .IN3(~na1191_2), .IN4(na1188_1), .IN5(~na1193_1), .IN6(1'b1), .IN7(~na1191_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x82y72     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7361_4 ( .OUT(na7361_2), .IN1(~na428_1), .IN2(1'b0), .IN3(~na9124_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y75     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7362_4 ( .OUT(na7362_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1530_1), .IN4(na2989_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x110y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7363_1 ( .OUT(na7363_1), .IN1(~na488_1), .IN2(~na1273_1), .IN3(~na8_2), .IN4(~na1210_1), .IN5(~na2667_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7364_1 ( .OUT(na7364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7364_6 ( .RAM_O1(na7364_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7364_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7365_4 ( .OUT(na7365_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7365_6 ( .RAM_O2(na7365_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7365_2), .COMP_OUT(1'b0) );
// C_AND////      x133y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7366_1 ( .OUT(na7366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7366_6 ( .RAM_O1(na7366_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7366_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x109y108     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7367_1 ( .OUT(na7367_1), .IN1(~na488_1), .IN2(~na1272_1), .IN3(~na8_2), .IN4(~na1209_1), .IN5(~na1109_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x133y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7368_4 ( .OUT(na7368_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7368_6 ( .RAM_O2(na7368_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7368_2), .COMP_OUT(1'b0) );
// C_AND////      x133y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7369_1 ( .OUT(na7369_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7369_6 ( .RAM_O1(na7369_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7369_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x128y35     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7370_2 ( .OUT(na7370_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6639_36), .CP_O(1'b0) );
// C_MX2b////      x61y124     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7371_1 ( .OUT(na7371_1), .IN1(na526_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1620_1), .IN6(na1393_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x108y101     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7372_1 ( .OUT(na7372_1), .IN1(~na488_1), .IN2(~na1271_1), .IN3(~na8_2), .IN4(~na1208_1), .IN5(~na1106_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x128y34     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7373_5 ( .OUT(na7373_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6639_37), .CP_O(1'b0) );
// C_/RAM_I1///      x128y34     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7374_2 ( .OUT(na7374_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6639_38), .CP_O(1'b0) );
// C_////RAM_I2      x128y33     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7375_5 ( .OUT(na7375_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6639_39), .CP_O(1'b0) );
// C_ORAND////      x104y104     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7376_1 ( .OUT(na7376_1), .IN1(~na488_1), .IN2(~na1269_1), .IN3(~na8_2), .IN4(~na1206_1), .IN5(~na1102_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x128y33     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7377_2 ( .OUT(na7377_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6639_40), .CP_O(1'b0) );
// C_AND////      x99y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7378_1 ( .OUT(na7378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7378_6 ( .RAM_O1(na7378_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7378_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y24     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7379_4 ( .OUT(na7379_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7379_6 ( .RAM_O2(na7379_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7379_2), .COMP_OUT(1'b0) );
// C_AND////      x92y24     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7380_1 ( .OUT(na7380_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7380_6 ( .RAM_O1(na7380_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7380_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x108y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7381_1 ( .OUT(na7381_1), .IN1(~na488_1), .IN2(~na1268_1), .IN3(~na8_2), .IN4(~na1205_1), .IN5(~na9650_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y23     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7382_4 ( .OUT(na7382_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7382_6 ( .RAM_O2(na7382_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7382_2), .COMP_OUT(1'b0) );
// C_AND////      x92y23     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7383_1 ( .OUT(na7383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7383_6 ( .RAM_O1(na7383_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7383_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y22     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7384_4 ( .OUT(na7384_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7384_6 ( .RAM_O2(na7384_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7384_2), .COMP_OUT(1'b0) );
// C_ORAND////      x102y101     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7385_1 ( .OUT(na7385_1), .IN1(~na488_1), .IN2(~na1267_1), .IN3(~na8_2), .IN4(~na1204_1), .IN5(~na1100_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y22     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7386_1 ( .OUT(na7386_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7386_6 ( .RAM_O1(na7386_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7386_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y21     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7387_4 ( .OUT(na7387_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7387_6 ( .RAM_O2(na7387_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7387_2), .COMP_OUT(1'b0) );
// C_AND////      x92y21     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7388_1 ( .OUT(na7388_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7388_6 ( .RAM_O1(na7388_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7388_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x104y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7389_1 ( .OUT(na7389_1), .IN1(~na488_1), .IN2(~na1266_1), .IN3(~na8_2), .IN4(~na1203_1), .IN5(~na1098_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y20     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7390_4 ( .OUT(na7390_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7390_6 ( .RAM_O2(na7390_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7390_2), .COMP_OUT(1'b0) );
// C_AND////      x92y20     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7391_1 ( .OUT(na7391_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7391_6 ( .RAM_O1(na7391_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7391_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y19     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7392_4 ( .OUT(na7392_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7392_6 ( .RAM_O2(na7392_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7392_2), .COMP_OUT(1'b0) );
// C_ORAND////      x106y99     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7393_1 ( .OUT(na7393_1), .IN1(~na488_1), .IN2(~na9480_2), .IN3(~na8_2), .IN4(~na9449_2), .IN5(~na9403_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y19     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7394_1 ( .OUT(na7394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7394_6 ( .RAM_O1(na7394_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7394_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y18     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7395_4 ( .OUT(na7395_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7395_6 ( .RAM_O2(na7395_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7395_2), .COMP_OUT(1'b0) );
// C_AND////      x92y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7396_1 ( .OUT(na7396_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7396_6 ( .RAM_O1(na7396_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7396_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x109y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7397_1 ( .OUT(na7397_1), .IN1(~na488_1), .IN2(~na1264_1), .IN3(~na8_2), .IN4(~na1201_1), .IN5(~na1094_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7398_4 ( .OUT(na7398_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7398_6 ( .RAM_O2(na7398_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7398_2), .COMP_OUT(1'b0) );
// C_AND////      x92y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7399_1 ( .OUT(na7399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7399_6 ( .RAM_O1(na7399_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7399_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y19     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7400_4 ( .OUT(na7400_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7400_6 ( .RAM_O2(na7400_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7400_2), .COMP_OUT(1'b0) );
// C_ORAND////      x106y100     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7401_1 ( .OUT(na7401_1), .IN1(~na488_1), .IN2(~na1263_1), .IN3(~na8_2), .IN4(~na1200_1), .IN5(~na1093_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y19     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7402_1 ( .OUT(na7402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7402_6 ( .RAM_O1(na7402_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7402_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7403_4 ( .OUT(na7403_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7403_6 ( .RAM_O2(na7403_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7403_2), .COMP_OUT(1'b0) );
// C_AND////      x101y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7404_1 ( .OUT(na7404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7404_6 ( .RAM_O1(na7404_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7404_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x110y101     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7405_1 ( .OUT(na7405_1), .IN1(~na488_1), .IN2(~na1262_1), .IN3(~na8_2), .IN4(~na1199_1), .IN5(~na1092_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7406_4 ( .OUT(na7406_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7406_6 ( .RAM_O2(na7406_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7406_2), .COMP_OUT(1'b0) );
// C_AND////      x101y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7407_1 ( .OUT(na7407_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7407_6 ( .RAM_O1(na7407_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7407_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x96y19     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7408_2 ( .OUT(na7408_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6640_36), .CP_O(1'b0) );
// C_ORAND////      x108y100     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7409_1 ( .OUT(na7409_1), .IN1(~na488_1), .IN2(~na1261_1), .IN3(~na8_2), .IN4(~na1198_1), .IN5(~na1090_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x96y18     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7410_5 ( .OUT(na7410_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6640_37), .CP_O(1'b0) );
// C_/RAM_I1///      x96y18     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7411_2 ( .OUT(na7411_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6640_38), .CP_O(1'b0) );
// C_////RAM_I2      x96y17     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7412_5 ( .OUT(na7412_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6640_39), .CP_O(1'b0) );
// C_ORAND////      x111y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7413_1 ( .OUT(na7413_1), .IN1(~na488_1), .IN2(~na1245_1), .IN3(~na8_2), .IN4(~na1197_1), .IN5(~na1089_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x96y17     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7414_2 ( .OUT(na7414_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6640_40), .CP_O(1'b0) );
// C_AND////      x35y113     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7415_1 ( .OUT(na7415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7415_6 ( .RAM_O1(na7415_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7415_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y120     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7416_4 ( .OUT(na7416_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7416_6 ( .RAM_O2(na7416_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7416_2), .COMP_OUT(1'b0) );
// C_ORAND////      x115y104     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7417_1 ( .OUT(na7417_1), .IN1(~na488_1), .IN2(~na1244_1), .IN3(~na8_2), .IN4(~na1164_1), .IN5(~na9400_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y120     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7418_1 ( .OUT(na7418_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7418_6 ( .RAM_O1(na7418_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7418_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y119     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7419_4 ( .OUT(na7419_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7419_6 ( .RAM_O2(na7419_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7419_2), .COMP_OUT(1'b0) );
// C_AND////      x28y119     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7420_1 ( .OUT(na7420_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7420_6 ( .RAM_O1(na7420_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7420_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x113y105     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7421_1 ( .OUT(na7421_1), .IN1(~na488_1), .IN2(~na1243_1), .IN3(~na8_2), .IN4(~na1163_1), .IN5(~na1087_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y118     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7422_4 ( .OUT(na7422_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7422_6 ( .RAM_O2(na7422_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7422_2), .COMP_OUT(1'b0) );
// C_AND////      x28y118     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7423_1 ( .OUT(na7423_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7423_6 ( .RAM_O1(na7423_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7423_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y117     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7424_4 ( .OUT(na7424_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7424_6 ( .RAM_O2(na7424_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7424_2), .COMP_OUT(1'b0) );
// C_ORAND////      x110y103     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7425_1 ( .OUT(na7425_1), .IN1(~na488_1), .IN2(~na1242_1), .IN3(~na8_2), .IN4(~na1162_1), .IN5(~na1086_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y117     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7426_1 ( .OUT(na7426_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7426_6 ( .RAM_O1(na7426_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7426_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y116     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7427_4 ( .OUT(na7427_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7427_6 ( .RAM_O2(na7427_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7427_2), .COMP_OUT(1'b0) );
// C_AND////      x28y116     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7428_1 ( .OUT(na7428_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7428_6 ( .RAM_O1(na7428_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7428_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x114y106     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7429_1 ( .OUT(na7429_1), .IN1(~na488_1), .IN2(~na1241_1), .IN3(~na8_2), .IN4(~na1161_1), .IN5(~na1081_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y115     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7430_4 ( .OUT(na7430_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7430_6 ( .RAM_O2(na7430_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7430_2), .COMP_OUT(1'b0) );
// C_AND////      x28y115     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7431_1 ( .OUT(na7431_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7431_6 ( .RAM_O1(na7431_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7431_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y114     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7432_4 ( .OUT(na7432_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7432_6 ( .RAM_O2(na7432_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7432_2), .COMP_OUT(1'b0) );
// C_ORAND////      x110y105     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7433_1 ( .OUT(na7433_1), .IN1(~na488_1), .IN2(~na1240_1), .IN3(~na8_2), .IN4(~na1159_1), .IN5(~na2669_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y114     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7434_1 ( .OUT(na7434_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7434_6 ( .RAM_O1(na7434_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7434_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y113     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7435_4 ( .OUT(na7435_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7435_6 ( .RAM_O2(na7435_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7435_2), .COMP_OUT(1'b0) );
// C_AND////      x28y113     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7436_1 ( .OUT(na7436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7436_6 ( .RAM_O1(na7436_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7436_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x112y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7437_1 ( .OUT(na7437_1), .IN1(~na488_1), .IN2(~na1238_1), .IN3(~na8_2), .IN4(~na1157_1), .IN5(~na1077_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y115     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7438_4 ( .OUT(na7438_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7438_6 ( .RAM_O2(na7438_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7438_2), .COMP_OUT(1'b0) );
// C_AND////      x37y115     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7439_1 ( .OUT(na7439_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7439_6 ( .RAM_O1(na7439_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7439_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y114     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7440_4 ( .OUT(na7440_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7440_6 ( .RAM_O2(na7440_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7440_2), .COMP_OUT(1'b0) );
// C_ORAND////      x113y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7441_1 ( .OUT(na7441_1), .IN1(~na488_1), .IN2(~na1239_1), .IN3(~na8_2), .IN4(~na9430_2), .IN5(~na1080_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y114     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7442_1 ( .OUT(na7442_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7442_6 ( .RAM_O1(na7442_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7442_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y113     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7443_4 ( .OUT(na7443_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7443_6 ( .RAM_O2(na7443_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7443_2), .COMP_OUT(1'b0) );
// C_AND////      x37y113     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7444_1 ( .OUT(na7444_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7444_6 ( .RAM_O1(na7444_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7444_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x114y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7445_1 ( .OUT(na7445_1), .IN1(~na488_1), .IN2(~na1234_1), .IN3(~na8_2), .IN4(~na1156_1), .IN5(~na1075_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x32y115     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7446_2 ( .OUT(na7446_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6641_36), .CP_O(1'b0) );
// C_////RAM_I2      x32y114     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7447_5 ( .OUT(na7447_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6641_37), .CP_O(1'b0) );
// C_/RAM_I1///      x32y114     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7448_2 ( .OUT(na7448_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6641_38), .CP_O(1'b0) );
// C_ORAND////      x114y107     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7449_1 ( .OUT(na7449_1), .IN1(~na488_1), .IN2(~na1233_1), .IN3(~na8_2), .IN4(~na1155_1), .IN5(~na9394_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x32y113     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7450_5 ( .OUT(na7450_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6641_39), .CP_O(1'b0) );
// C_/RAM_I1///      x32y113     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7451_2 ( .OUT(na7451_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6641_40), .CP_O(1'b0) );
// C_AND////      x35y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7452_1 ( .OUT(na7452_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7452_6 ( .RAM_O1(na7452_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7452_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x115y106     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7453_1 ( .OUT(na7453_1), .IN1(~na488_1), .IN2(~na1232_1), .IN3(~na8_2), .IN4(~na9424_2), .IN5(~na1072_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y24     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7454_4 ( .OUT(na7454_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7454_6 ( .RAM_O2(na7454_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7454_2), .COMP_OUT(1'b0) );
// C_AND////      x28y24     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7455_1 ( .OUT(na7455_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7455_6 ( .RAM_O1(na7455_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7455_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y23     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7456_4 ( .OUT(na7456_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7456_6 ( .RAM_O2(na7456_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7456_2), .COMP_OUT(1'b0) );
// C_ORAND////      x110y100     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7457_1 ( .OUT(na7457_1), .IN1(~na488_1), .IN2(~na1231_1), .IN3(~na8_2), .IN4(~na9422_2), .IN5(~na1071_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y23     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7458_1 ( .OUT(na7458_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7458_6 ( .RAM_O1(na7458_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7458_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y22     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7459_4 ( .OUT(na7459_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7459_6 ( .RAM_O2(na7459_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7459_2), .COMP_OUT(1'b0) );
// C_AND////      x28y22     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7460_1 ( .OUT(na7460_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7460_6 ( .RAM_O1(na7460_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7460_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x102y105     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7461_1 ( .OUT(na7461_1), .IN1(~na488_1), .IN2(~na1230_1), .IN3(~na8_2), .IN4(~na1152_1), .IN5(~na1070_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y21     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7462_4 ( .OUT(na7462_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7462_6 ( .RAM_O2(na7462_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7462_2), .COMP_OUT(1'b0) );
// C_AND////      x28y21     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7463_1 ( .OUT(na7463_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7463_6 ( .RAM_O1(na7463_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7463_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y20     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7464_4 ( .OUT(na7464_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7464_6 ( .RAM_O2(na7464_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7464_2), .COMP_OUT(1'b0) );
// C_ORAND////      x113y96     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7465_1 ( .OUT(na7465_1), .IN1(~na488_1), .IN2(~na1229_1), .IN3(~na8_2), .IN4(~na1151_1), .IN5(~na1069_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y20     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7466_1 ( .OUT(na7466_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7466_6 ( .RAM_O1(na7466_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7466_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y19     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7467_4 ( .OUT(na7467_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7467_6 ( .RAM_O2(na7467_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7467_2), .COMP_OUT(1'b0) );
// C_AND////      x28y19     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7468_1 ( .OUT(na7468_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7468_6 ( .RAM_O1(na7468_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7468_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x111y98     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7469_1 ( .OUT(na7469_1), .IN1(~na488_1), .IN2(~na1228_1), .IN3(~na8_2), .IN4(~na1150_1), .IN5(~na1068_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y18     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7470_4 ( .OUT(na7470_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7470_6 ( .RAM_O2(na7470_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7470_2), .COMP_OUT(1'b0) );
// C_AND////      x28y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7471_1 ( .OUT(na7471_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7471_6 ( .RAM_O1(na7471_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7471_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7472_4 ( .OUT(na7472_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7472_6 ( .RAM_O2(na7472_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7472_2), .COMP_OUT(1'b0) );
// C_ORAND////      x110y98     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7473_1 ( .OUT(na7473_1), .IN1(~na488_1), .IN2(~na1227_1), .IN3(~na8_2), .IN4(~na1149_1), .IN5(~na2670_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7474_1 ( .OUT(na7474_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7474_6 ( .RAM_O1(na7474_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7474_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y19     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7475_4 ( .OUT(na7475_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7475_6 ( .RAM_O2(na7475_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7475_2), .COMP_OUT(1'b0) );
// C_AND////      x37y19     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7476_1 ( .OUT(na7476_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7476_6 ( .RAM_O1(na7476_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7476_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x110y97     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7477_1 ( .OUT(na7477_1), .IN1(~na488_1), .IN2(~na1226_1), .IN3(~na8_2), .IN4(~na1148_1), .IN5(~na1035_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7478_4 ( .OUT(na7478_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7478_6 ( .RAM_O2(na7478_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7478_2), .COMP_OUT(1'b0) );
// C_AND////      x37y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7479_1 ( .OUT(na7479_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7479_6 ( .RAM_O1(na7479_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7479_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7480_4 ( .OUT(na7480_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7480_6 ( .RAM_O2(na7480_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7480_2), .COMP_OUT(1'b0) );
// C_ORAND////      x108y98     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7481_1 ( .OUT(na7481_1), .IN1(~na488_1), .IN2(~na2666_1), .IN3(~na8_2), .IN4(~na1147_1), .IN5(~na1032_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7482_1 ( .OUT(na7482_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7482_6 ( .RAM_O1(na7482_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7482_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x32y19     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7483_2 ( .OUT(na7483_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6642_36), .CP_O(1'b0) );
// C_////RAM_I2      x32y18     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7484_5 ( .OUT(na7484_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6642_37), .CP_O(1'b0) );
// C_OR////      x86y89     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7485_1 ( .OUT(na7485_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1145_1), .IN8(~na1531_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y85     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7486_4 ( .OUT(na7486_2), .IN1(1'b1), .IN2(na1595_2), .IN3(na1213_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x87y89     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7487_4 ( .OUT(na7487_2), .IN1(~na1274_1), .IN2(~na1612_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y73     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7488_4 ( .OUT(na7488_2), .IN1(na1028_1), .IN2(1'b1), .IN3(na1026_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y100     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7489_1 ( .OUT(na7489_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na428_1), .IN6(1'b0), .IN7(~na1030_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y96     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7490_4 ( .OUT(na7490_2), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1527_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x92y92     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7491_1 ( .OUT(na7491_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1216_1), .IN6(1'b0), .IN7(~na1530_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y100     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7492_4 ( .OUT(na7492_2), .IN1(1'b1), .IN2(na1524_1), .IN3(na1275_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y83     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7493_1 ( .OUT(na7493_1), .IN1(~na488_1), .IN2(~na3109_1), .IN3(~na8_2), .IN4(~na3017_1), .IN5(~na3001_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x32y18     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7494_2 ( .OUT(na7494_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6642_38), .CP_O(1'b0) );
// C_////RAM_I2      x32y17     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7495_5 ( .OUT(na7495_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6642_39), .CP_O(1'b0) );
// C_/RAM_I1///      x32y17     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7496_2 ( .OUT(na7496_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6642_40), .CP_O(1'b0) );
// C_ORAND////      x108y95     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7497_1 ( .OUT(na7497_1), .IN1(~na488_1), .IN2(~na3111_1), .IN3(~na8_2), .IN4(~na3071_1), .IN5(~na990_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x131y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7498_1 ( .OUT(na7498_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7498_6 ( .RAM_O1(na7498_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7498_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y24     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7499_4 ( .OUT(na7499_2), .IN1(1'b1), .IN2(1'b1), .IN3(na90_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7499_6 ( .RAM_O2(na7499_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7499_2), .COMP_OUT(1'b0) );
// C_AND////      x124y24     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7500_1 ( .OUT(na7500_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7500_6 ( .RAM_O1(na7500_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7500_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x120y89     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7501_1 ( .OUT(na7501_1), .IN1(~na488_1), .IN2(~na3112_1), .IN3(~na8_2), .IN4(~na3072_1), .IN5(~na1883_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y23     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7502_4 ( .OUT(na7502_2), .IN1(na88_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7502_6 ( .RAM_O2(na7502_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7502_2), .COMP_OUT(1'b0) );
// C_AND////      x124y23     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7503_1 ( .OUT(na7503_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7503_6 ( .RAM_O1(na7503_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7503_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y22     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7504_4 ( .OUT(na7504_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7504_6 ( .RAM_O2(na7504_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7504_2), .COMP_OUT(1'b0) );
// C_ORAND////      x99y83     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7505_1 ( .OUT(na7505_1), .IN1(~na488_1), .IN2(~na570_1), .IN3(~na8_2), .IN4(~na3073_1), .IN5(~na1868_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y22     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7506_1 ( .OUT(na7506_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7506_6 ( .RAM_O1(na7506_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7506_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y21     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7507_4 ( .OUT(na7507_2), .IN1(1'b1), .IN2(1'b1), .IN3(na84_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7507_6 ( .RAM_O2(na7507_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7507_2), .COMP_OUT(1'b0) );
// C_AND////      x124y21     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7508_1 ( .OUT(na7508_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7508_6 ( .RAM_O1(na7508_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7508_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x110y77     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7509_1 ( .OUT(na7509_1), .IN1(~na488_1), .IN2(~na639_1), .IN3(~na8_2), .IN4(~na3074_1), .IN5(~na1138_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y20     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7510_4 ( .OUT(na7510_2), .IN1(1'b1), .IN2(na35_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7510_6 ( .RAM_O2(na7510_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7510_2), .COMP_OUT(1'b0) );
// C_AND////      x124y20     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7511_1 ( .OUT(na7511_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na37_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7511_6 ( .RAM_O1(na7511_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7511_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y19     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7512_4 ( .OUT(na7512_2), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7512_6 ( .RAM_O2(na7512_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7512_2), .COMP_OUT(1'b0) );
// C_ORAND////      x116y88     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7513_1 ( .OUT(na7513_1), .IN1(~na488_1), .IN2(~na785_1), .IN3(~na8_2), .IN4(~na3075_1), .IN5(~na1869_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y19     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7514_1 ( .OUT(na7514_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na66_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7514_6 ( .RAM_O1(na7514_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7514_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x124y18     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7515_4 ( .OUT(na7515_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7515_6 ( .RAM_O2(na7515_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7515_2), .COMP_OUT(1'b0) );
// C_AND////      x124y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7516_1 ( .OUT(na7516_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7516_6 ( .RAM_O1(na7516_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7516_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x115y79     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7517_1 ( .OUT(na7517_1), .IN1(~na488_1), .IN2(~na827_1), .IN3(~na8_2), .IN4(~na3076_1), .IN5(~na2906_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x124y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7518_4 ( .OUT(na7518_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7518_6 ( .RAM_O2(na7518_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7518_2), .COMP_OUT(1'b0) );
// C_AND////      x124y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7519_1 ( .OUT(na7519_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7519_6 ( .RAM_O1(na7519_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7519_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y19     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7520_4 ( .OUT(na7520_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7520_6 ( .RAM_O2(na7520_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7520_2), .COMP_OUT(1'b0) );
// C_ORAND////      x113y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7521_1 ( .OUT(na7521_1), .IN1(~na488_1), .IN2(~na1371_1), .IN3(~na8_2), .IN4(~na9754_2), .IN5(~na3212_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x133y19     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7522_1 ( .OUT(na7522_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7522_6 ( .RAM_O1(na7522_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7522_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x133y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7523_4 ( .OUT(na7523_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7523_6 ( .RAM_O2(na7523_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7523_2), .COMP_OUT(1'b0) );
// C_AND////      x133y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7524_1 ( .OUT(na7524_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7524_6 ( .RAM_O1(na7524_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7524_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x114y81     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7525_1 ( .OUT(na7525_1), .IN1(~na488_1), .IN2(~na1411_1), .IN3(~na8_2), .IN4(~na3117_1), .IN5(~na2246_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x133y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7526_4 ( .OUT(na7526_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7526_6 ( .RAM_O2(na7526_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7526_2), .COMP_OUT(1'b0) );
// C_AND////      x133y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7527_1 ( .OUT(na7527_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7527_6 ( .RAM_O1(na7527_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7527_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x128y19     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7528_2 ( .OUT(na7528_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6643_36), .CP_O(1'b0) );
// C_ORAND////      x117y83     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7529_1 ( .OUT(na7529_1), .IN1(~na488_1), .IN2(~na1693_1), .IN3(~na8_2), .IN4(~na3123_1), .IN5(~na2254_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x128y18     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7530_5 ( .OUT(na7530_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6643_37), .CP_O(1'b0) );
// C_/RAM_I1///      x128y18     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7531_2 ( .OUT(na7531_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6643_38), .CP_O(1'b0) );
// C_////RAM_I2      x128y17     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7532_5 ( .OUT(na7532_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6643_39), .CP_O(1'b0) );
// C_ORAND////      x116y83     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7533_1 ( .OUT(na7533_1), .IN1(~na488_1), .IN2(~na9706_2), .IN3(~na8_2), .IN4(~na9759_2), .IN5(~na2717_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x128y17     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a7534_2 ( .OUT(na7534_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6643_40), .CP_O(1'b0) );
// C_AND////      x67y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7535_1 ( .OUT(na7535_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7535_6 ( .RAM_O1(na7535_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7535_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x59y97     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7536_4 ( .OUT(na7536_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3273_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7536_6 ( .RAM_O2(na7536_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7536_2), .COMP_OUT(1'b0) );
// C_ORAND////      x114y95     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7537_1 ( .OUT(na7537_1), .IN1(~na488_1), .IN2(~na2909_1), .IN3(~na8_2), .IN4(~na9762_2), .IN5(~na2745_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y104     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7538_4 ( .OUT(na7538_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7538_6 ( .RAM_O2(na7538_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7538_2), .COMP_OUT(1'b0) );
// C_AND////      x60y104     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7539_1 ( .OUT(na7539_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7539_6 ( .RAM_O1(na7539_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7539_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y103     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7540_4 ( .OUT(na7540_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7540_6 ( .RAM_O2(na7540_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7540_2), .COMP_OUT(1'b0) );
// C_ORAND////      x112y87     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7541_1 ( .OUT(na7541_1), .IN1(~na488_1), .IN2(~na2910_1), .IN3(~na8_2), .IN4(~na3129_1), .IN5(~na471_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y103     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7542_1 ( .OUT(na7542_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7542_6 ( .RAM_O1(na7542_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7542_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y102     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7543_4 ( .OUT(na7543_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7543_6 ( .RAM_O2(na7543_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7543_2), .COMP_OUT(1'b0) );
// C_AND////      x60y102     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7544_1 ( .OUT(na7544_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7544_6 ( .RAM_O1(na7544_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7544_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x121y85     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7545_1 ( .OUT(na7545_1), .IN1(~na488_1), .IN2(~na2911_1), .IN3(~na8_2), .IN4(~na579_1), .IN5(~na1726_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y101     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7546_4 ( .OUT(na7546_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7546_6 ( .RAM_O2(na7546_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7546_2), .COMP_OUT(1'b0) );
// C_AND////      x60y101     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7547_1 ( .OUT(na7547_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7547_6 ( .RAM_O1(na7547_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7547_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y100     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7548_4 ( .OUT(na7548_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7548_6 ( .RAM_O2(na7548_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7548_2), .COMP_OUT(1'b0) );
// C_ORAND////      x119y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7549_1 ( .OUT(na7549_1), .IN1(~na488_1), .IN2(~na9709_2), .IN3(~na8_2), .IN4(~na663_1), .IN5(~na457_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y100     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7550_1 ( .OUT(na7550_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7550_6 ( .RAM_O1(na7550_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7550_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y99     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7551_4 ( .OUT(na7551_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7551_6 ( .RAM_O2(na7551_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7551_2), .COMP_OUT(1'b0) );
// C_AND////      x60y99     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7552_1 ( .OUT(na7552_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7552_6 ( .RAM_O1(na7552_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7552_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x122y85     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7553_1 ( .OUT(na7553_1), .IN1(~na488_1), .IN2(~na9710_2), .IN3(~na8_2), .IN4(~na9336_2), .IN5(~na3211_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y98     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7554_4 ( .OUT(na7554_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7554_6 ( .RAM_O2(na7554_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7554_2), .COMP_OUT(1'b0) );
// C_AND////      x60y98     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7555_1 ( .OUT(na7555_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7555_6 ( .RAM_O1(na7555_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7555_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y97     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7556_4 ( .OUT(na7556_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7556_6 ( .RAM_O2(na7556_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7556_2), .COMP_OUT(1'b0) );
// C_ORAND////      x114y85     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7557_1 ( .OUT(na7557_1), .IN1(~na488_1), .IN2(~na2936_1), .IN3(~na8_2), .IN4(~na1512_1), .IN5(~na3193_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7558_1 ( .OUT(na7558_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7558_6 ( .RAM_O1(na7558_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7558_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y100     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7559_1 ( .OUT(na7559_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7559_6 ( .RAM_O1(na7559_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7559_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y99     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7560_1 ( .OUT(na7560_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7560_6 ( .RAM_O1(na7560_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7560_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x123y83     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7561_1 ( .OUT(na7561_1), .IN1(~na488_1), .IN2(~na9716_2), .IN3(~na8_2), .IN4(~na9673_2), .IN5(~na3171_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y98     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7562_4 ( .OUT(na7562_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7562_6 ( .RAM_O2(na7562_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7562_2), .COMP_OUT(1'b0) );
// C_AND////      x69y98     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7563_1 ( .OUT(na7563_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7563_6 ( .RAM_O1(na7563_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7563_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y97     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7564_4 ( .OUT(na7564_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7564_6 ( .RAM_O2(na7564_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7564_2), .COMP_OUT(1'b0) );
// C_ORAND////      x117y86     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7565_1 ( .OUT(na7565_1), .IN1(~na488_1), .IN2(~na2944_1), .IN3(~na8_2), .IN4(~na2661_1), .IN5(~na3166_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y97     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7566_1 ( .OUT(na7566_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7566_6 ( .RAM_O1(na7566_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7566_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y104     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7567_4 ( .OUT(na7567_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7567_5 ( .OUT(na7567_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7567_6 ( .RAM_O2(na7567_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7567_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y104     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7568_1 ( .OUT(na7568_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7568_2 ( .OUT(na7568_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7568_6 ( .RAM_O1(na7568_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7568_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x112y97     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7569_1 ( .OUT(na7569_1), .IN1(~na488_1), .IN2(~na2945_1), .IN3(~na8_2), .IN4(~na3189_1), .IN5(~na9770_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x62y103     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7570_4 ( .OUT(na7570_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7570_5 ( .OUT(na7570_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7570_6 ( .RAM_O2(na7570_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7570_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y103     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7571_1 ( .OUT(na7571_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7571_2 ( .OUT(na7571_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7571_6 ( .RAM_O1(na7571_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7571_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y104     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7572_4 ( .OUT(na7572_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7572_5 ( .OUT(na7572_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7572_6 ( .RAM_O2(na7572_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7572_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x110y87     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7573_1 ( .OUT(na7573_1), .IN1(~na488_1), .IN2(~na2946_1), .IN3(~na8_2), .IN4(~na9785_2), .IN5(~na3150_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y104     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7574_1 ( .OUT(na7574_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7574_2 ( .OUT(na7574_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7574_6 ( .RAM_O1(na7574_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7574_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y103     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7575_4 ( .OUT(na7575_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7575_5 ( .OUT(na7575_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7575_6 ( .RAM_O2(na7575_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7575_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y103     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7576_1 ( .OUT(na7576_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7576_2 ( .OUT(na7576_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7576_6 ( .RAM_O1(na7576_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7576_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x116y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7577_1 ( .OUT(na7577_1), .IN1(~na488_1), .IN2(~na2955_1), .IN3(~na8_2), .IN4(~na3175_1), .IN5(~na2156_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y102     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7578_4 ( .OUT(na7578_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7578_5 ( .OUT(na7578_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7578_6 ( .RAM_O2(na7578_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7578_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y102     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7579_1 ( .OUT(na7579_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7579_2 ( .OUT(na7579_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7579_6 ( .RAM_O1(na7579_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7579_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y101     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7580_4 ( .OUT(na7580_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7580_5 ( .OUT(na7580_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7580_6 ( .RAM_O2(na7580_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7580_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x116y85     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7581_1 ( .OUT(na7581_1), .IN1(~na488_1), .IN2(~na2956_1), .IN3(~na8_2), .IN4(~na3165_1), .IN5(~na1889_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y101     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7582_1 ( .OUT(na7582_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7582_2 ( .OUT(na7582_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7582_6 ( .RAM_O1(na7582_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7582_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y100     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7583_4 ( .OUT(na7583_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7583_5 ( .OUT(na7583_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7583_6 ( .RAM_O2(na7583_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7583_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y100     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7584_1 ( .OUT(na7584_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7584_2 ( .OUT(na7584_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7584_6 ( .RAM_O1(na7584_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7584_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x114y87     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7585_1 ( .OUT(na7585_1), .IN1(~na488_1), .IN2(~na2957_1), .IN3(~na8_2), .IN4(~na3156_1), .IN5(~na3136_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y99     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7586_4 ( .OUT(na7586_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7586_5 ( .OUT(na7586_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7586_6 ( .RAM_O2(na7586_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7586_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y99     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7587_1 ( .OUT(na7587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7587_2 ( .OUT(na7587_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7587_6 ( .RAM_O1(na7587_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7587_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y98     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7588_4 ( .OUT(na7588_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7588_5 ( .OUT(na7588_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7588_6 ( .RAM_O2(na7588_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7588_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x110y79     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7589_1 ( .OUT(na7589_1), .IN1(~na488_1), .IN2(~na9733_2), .IN3(~na8_2), .IN4(~na9774_2), .IN5(~na1697_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y98     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7590_1 ( .OUT(na7590_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7590_2 ( .OUT(na7590_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7590_6 ( .RAM_O1(na7590_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7590_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y97     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7591_4 ( .OUT(na7591_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7591_5 ( .OUT(na7591_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7591_6 ( .RAM_O2(na7591_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7591_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y97     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7592_1 ( .OUT(na7592_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7592_2 ( .OUT(na7592_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6644_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7592_6 ( .RAM_O1(na7592_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7592_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x96y80     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7593_1 ( .OUT(na7593_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1891_1), .IN8(~na1531_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y84     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7594_4 ( .OUT(na7594_2), .IN1(1'b1), .IN2(na1595_2), .IN3(na3014_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y83     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7595_1 ( .OUT(na7595_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1612_1), .IN7(1'b0), .IN8(~na9750_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y61     80'h00_0018_00_0000_0888_F42A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7596_1 ( .OUT(na7596_1), .IN1(na1045_2), .IN2(1'b1), .IN3(na3186_2), .IN4(~na37_1), .IN5(~na86_1), .IN6(na69_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x99y84     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7597_4 ( .OUT(na7597_2), .IN1(~na428_1), .IN2(1'b0), .IN3(~na1892_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y84     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7598_1 ( .OUT(na7598_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3178_2), .IN7(1'b1), .IN8(na1527_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x98y77     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7599_1 ( .OUT(na7599_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3012_1), .IN6(1'b0), .IN7(~na1530_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x102y69     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7600_4 ( .OUT(na7600_2), .IN1(1'b1), .IN2(na1524_1), .IN3(na9510_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y106     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7601_1 ( .OUT(na7601_1), .IN1(~na853_2), .IN2(~na9356_2), .IN3(~na8_2), .IN4(~na4907_2), .IN5(~na9357_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y104     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7602_4 ( .OUT(na7602_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2846_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7602_6 ( .RAM_O2(na7602_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7602_2), .COMP_OUT(1'b0) );
// C_AND////      x61y104     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7603_1 ( .OUT(na7603_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2846_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7603_6 ( .RAM_O1(na7603_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7603_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y103     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7604_4 ( .OUT(na7604_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2846_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7604_6 ( .RAM_O2(na7604_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7604_2), .COMP_OUT(1'b0) );
// C_ORAND////      x91y108     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7605_1 ( .OUT(na7605_1), .IN1(~na853_2), .IN2(~na9353_2), .IN3(~na8_2), .IN4(~na4905_2), .IN5(~na9354_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x61y103     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7606_1 ( .OUT(na7606_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2846_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7606_6 ( .RAM_O1(na7606_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7606_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y104     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7607_4 ( .OUT(na7607_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2844_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7607_6 ( .RAM_O2(na7607_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7607_2), .COMP_OUT(1'b0) );
// C_AND////      x63y104     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7608_1 ( .OUT(na7608_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2844_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7608_6 ( .RAM_O1(na7608_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7608_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x115y71     80'h00_0018_00_0000_0CEE_0700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7609_1 ( .OUT(na7609_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2825_1), .IN6(~na1042_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x125y72     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7610_4 ( .OUT(na7610_2), .IN1(1'b1), .IN2(1'b1), .IN3(na8_2), .IN4(na6095_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x117y72     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7611_1 ( .OUT(na7611_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na2824_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x123y71     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7612_4 ( .OUT(na7612_2), .IN1(1'b1), .IN2(1'b1), .IN3(na8_2), .IN4(na6096_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x115y70     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7613_4 ( .OUT(na7613_2), .IN1(1'b0), .IN2(~na1042_1), .IN3(1'b0), .IN4(~na2826_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x119y69     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7614_1 ( .OUT(na7614_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na6094_1), .IN6(1'b1), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x113y70     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7615_1 ( .OUT(na7615_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na2823_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x119y73     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7616_1 ( .OUT(na7616_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6097_2), .IN7(na8_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x113y64     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7617_1 ( .OUT(na7617_1), .IN1(~na2832_1), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na6093_2), .IN5(~na9693_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y103     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7618_4 ( .OUT(na7618_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2844_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7618_6 ( .RAM_O2(na7618_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7618_2), .COMP_OUT(1'b0) );
// C_AND////      x63y103     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7619_1 ( .OUT(na7619_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2844_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7619_6 ( .RAM_O1(na7619_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7619_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y102     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7620_4 ( .OUT(na7620_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2844_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7620_6 ( .RAM_O2(na7620_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7620_2), .COMP_OUT(1'b0) );
// C_///OR/      x105y72     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7621_4 ( .OUT(na7621_2), .IN1(~na2821_1), .IN2(~na1042_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x121y77     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7622_1 ( .OUT(na7622_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na8_2), .IN8(na6098_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x109y64     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7623_1 ( .OUT(na7623_1), .IN1(~na2833_1), .IN2(~na955_1), .IN3(~na8_2), .IN4(~na6092_1), .IN5(~na2828_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x63y102     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7624_1 ( .OUT(na7624_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2844_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7624_6 ( .RAM_O1(na7624_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7624_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y101     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7625_4 ( .OUT(na7625_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2844_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7625_6 ( .RAM_O2(na7625_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7625_2), .COMP_OUT(1'b0) );
// C_AND////      x63y101     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7626_1 ( .OUT(na7626_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2844_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7626_6 ( .RAM_O1(na7626_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7626_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x114y65     80'h00_0018_00_0000_0888_1C5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7627_1 ( .OUT(na7627_1), .IN1(1'b1), .IN2(na7629_2), .IN3(~na7628_2), .IN4(1'b1), .IN5(1'b1), .IN6(na7629_1), .IN7(~na7632_2),
                      .IN8(~na7630_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y73     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7628_4 ( .OUT(na7628_2), .IN1(na853_2), .IN2(na2760_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x119y68     80'h00_0078_00_0000_0CEE_3353
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7629_1 ( .OUT(na7629_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1042_1), .IN7(1'b0), .IN8(~na2829_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7629_4 ( .OUT(na7629_2), .IN1(1'b0), .IN2(~na6091_2), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y74     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7630_1 ( .OUT(na7630_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na488_1), .IN6(1'b1), .IN7(na2830_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y100     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7631_4 ( .OUT(na7631_2), .IN1(na2839_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7631_6 ( .RAM_O2(na7631_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7631_2), .COMP_OUT(1'b0) );
// C_///AND/      x120y61     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7632_4 ( .OUT(na7632_2), .IN1(1'b1), .IN2(na2834_1), .IN3(1'b1), .IN4(na9362_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y103     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7633_1 ( .OUT(na7633_1), .IN1(~na853_2), .IN2(~na9488_2), .IN3(~na8_2), .IN4(~na4903_2), .IN5(~na9489_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x63y100     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7634_1 ( .OUT(na7634_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2839_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7634_6 ( .RAM_O1(na7634_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7634_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y99     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7635_4 ( .OUT(na7635_2), .IN1(na2839_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7635_6 ( .RAM_O2(na7635_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7635_2), .COMP_OUT(1'b0) );
// C_AND////      x63y99     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7636_1 ( .OUT(na7636_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2839_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7636_6 ( .RAM_O1(na7636_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7636_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x92y107     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7637_1 ( .OUT(na7637_1), .IN1(~na853_2), .IN2(~na9655_2), .IN3(~na8_2), .IN4(~na4895_2), .IN5(~na9656_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y98     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7638_4 ( .OUT(na7638_2), .IN1(na2839_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7638_6 ( .RAM_O2(na7638_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7638_2), .COMP_OUT(1'b0) );
// C_AND////      x63y98     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7639_1 ( .OUT(na7639_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2839_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7639_6 ( .RAM_O1(na7639_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7639_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y97     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7640_4 ( .OUT(na7640_2), .IN1(na2839_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7640_6 ( .RAM_O2(na7640_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7640_2), .COMP_OUT(1'b0) );
// C_ORAND////      x84y80     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7641_1 ( .OUT(na7641_1), .IN1(~na853_2), .IN2(~na9495_2), .IN3(~na8_2), .IN4(~na4915_2), .IN5(~na9496_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x63y97     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7642_1 ( .OUT(na7642_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2839_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7642_6 ( .RAM_O1(na7642_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7642_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x99y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7643_1 ( .OUT(na7643_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7643_6 ( .RAM_O1(na7643_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7643_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x99y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7644_1 ( .OUT(na7644_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7644_6 ( .RAM_O1(na7644_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7644_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x90y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7645_1 ( .OUT(na7645_1), .IN1(~na853_2), .IN2(~na9497_2), .IN3(~na8_2), .IN4(~na4913_2), .IN5(~na9498_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y41     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7646_4 ( .OUT(na7646_2), .IN1(1'b1), .IN2(na3247_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7646_6 ( .RAM_O2(na7646_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7646_2), .COMP_OUT(1'b0) );
// C_///AND/      x91y33     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7647_4 ( .OUT(na7647_2), .IN1(1'b1), .IN2(na3249_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7647_6 ( .RAM_O2(na7647_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7647_2), .COMP_OUT(1'b0) );
// C_///AND/      x92y40     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7648_4 ( .OUT(na7648_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7648_6 ( .RAM_O2(na7648_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7648_2), .COMP_OUT(1'b0) );
// C_ORAND////      x86y84     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7649_1 ( .OUT(na7649_1), .IN1(~na853_2), .IN2(~na9657_2), .IN3(~na8_2), .IN4(~na4911_2), .IN5(~na9658_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y40     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7650_1 ( .OUT(na7650_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7650_6 ( .RAM_O1(na7650_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7650_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y39     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7651_4 ( .OUT(na7651_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7651_6 ( .RAM_O2(na7651_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7651_2), .COMP_OUT(1'b0) );
// C_AND////      x92y39     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7652_1 ( .OUT(na7652_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7652_6 ( .RAM_O1(na7652_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7652_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x87y85     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7653_1 ( .OUT(na7653_1), .IN1(~na853_2), .IN2(~na9390_2), .IN3(~na8_2), .IN4(~na4909_2), .IN5(~na9391_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y38     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7654_4 ( .OUT(na7654_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7654_6 ( .RAM_O2(na7654_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7654_2), .COMP_OUT(1'b0) );
// C_AND////      x92y38     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7655_1 ( .OUT(na7655_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7655_6 ( .RAM_O1(na7655_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7655_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y37     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7656_4 ( .OUT(na7656_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7656_6 ( .RAM_O2(na7656_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7656_2), .COMP_OUT(1'b0) );
// C_ORAND////      x91y105     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7657_1 ( .OUT(na7657_1), .IN1(~na853_2), .IN2(~na9385_2), .IN3(~na8_2), .IN4(~na4877_2), .IN5(~na9386_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y37     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7658_1 ( .OUT(na7658_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7658_6 ( .RAM_O1(na7658_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7658_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y36     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7659_4 ( .OUT(na7659_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7659_6 ( .RAM_O2(na7659_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7659_2), .COMP_OUT(1'b0) );
// C_AND////      x92y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7660_1 ( .OUT(na7660_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7660_6 ( .RAM_O1(na7660_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7660_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x105y93     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7661_1 ( .OUT(na7661_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3174_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y98     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7662_4 ( .OUT(na7662_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2255_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x105y96     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7663_4 ( .OUT(na7663_2), .IN1(~na3158_1), .IN2(1'b0), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y101     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7664_4 ( .OUT(na7664_2), .IN1(na853_2), .IN2(1'b1), .IN3(na2748_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x107y92     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7665_1 ( .OUT(na7665_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3132_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y97     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7666_4 ( .OUT(na7666_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na322_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x107y95     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7667_1 ( .OUT(na7667_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2797_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y110     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7668_4 ( .OUT(na7668_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2739_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y102     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7669_1 ( .OUT(na7669_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na2165_1), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y107     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7670_4 ( .OUT(na7670_2), .IN1(na853_2), .IN2(1'b1), .IN3(na247_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x103y98     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7671_1 ( .OUT(na7671_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1803_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y109     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7672_1 ( .OUT(na7672_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(na3205_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y92     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7673_1 ( .OUT(na7673_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1124_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y103     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7674_4 ( .OUT(na7674_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3201_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y89     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7675_1 ( .OUT(na7675_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na992_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y108     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7676_4 ( .OUT(na7676_2), .IN1(na853_2), .IN2(1'b1), .IN3(na3147_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x101y100     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7677_1 ( .OUT(na7677_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na960_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y107     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7678_4 ( .OUT(na7678_2), .IN1(na1903_1), .IN2(1'b1), .IN3(na9344_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y94     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7679_1 ( .OUT(na7679_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1867_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y107     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7680_4 ( .OUT(na7680_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3139_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x97y98     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7681_1 ( .OUT(na7681_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na558_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y105     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7682_4 ( .OUT(na7682_2), .IN1(na853_2), .IN2(1'b1), .IN3(na3134_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x109y96     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7683_1 ( .OUT(na7683_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na890_1), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y125     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7684_4 ( .OUT(na7684_2), .IN1(na1695_1), .IN2(na9345_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x107y94     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7685_1 ( .OUT(na7685_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na483_1), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y123     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7686_4 ( .OUT(na7686_2), .IN1(na853_2), .IN2(na3126_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y99     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7687_1 ( .OUT(na7687_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2720_1), .IN6(1'b0), .IN7(~na8_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y108     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7688_1 ( .OUT(na7688_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(na1656_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x105y97     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7689_4 ( .OUT(na7689_2), .IN1(~na2744_1), .IN2(1'b0), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y106     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7690_4 ( .OUT(na7690_2), .IN1(na853_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3130_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x115y103     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7691_4 ( .OUT(na7691_2), .IN1(~na447_1), .IN2(1'b0), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y104     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7692_1 ( .OUT(na7692_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(1'b1), .IN7(na1829_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x105y99     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7693_4 ( .OUT(na7693_2), .IN1(1'b0), .IN2(~na2251_1), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y108     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7694_1 ( .OUT(na7694_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(na3138_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x107y103     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7695_4 ( .OUT(na7695_2), .IN1(~na2170_1), .IN2(1'b0), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y108     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7696_1 ( .OUT(na7696_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(1'b1), .IN7(na3141_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x103y89     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7697_4 ( .OUT(na7697_2), .IN1(~na3210_1), .IN2(1'b0), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y106     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7698_1 ( .OUT(na7698_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3146_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x111y93     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7699_1 ( .OUT(na7699_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na8_2), .IN8(~na3207_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y106     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7700_1 ( .OUT(na7700_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(na3148_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x101y96     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7701_4 ( .OUT(na7701_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na8_2), .IN4(~na3197_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y107     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7702_1 ( .OUT(na7702_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(1'b1), .IN7(na2157_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x107y89     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7703_4 ( .OUT(na7703_2), .IN1(~na3194_1), .IN2(1'b0), .IN3(~na8_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y110     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7704_1 ( .OUT(na7704_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3169_1), .IN6(1'b1), .IN7(na9344_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x105y89     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7705_4 ( .OUT(na7705_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na8_2), .IN4(~na3172_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y106     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7706_1 ( .OUT(na7706_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na853_2), .IN6(1'b1), .IN7(na3190_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x109y87     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7707_4 ( .OUT(na7707_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na8_2), .IN4(~na3168_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y100     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7708_4 ( .OUT(na7708_2), .IN1(na853_2), .IN2(1'b1), .IN3(na3195_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x94y106     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7709_1 ( .OUT(na7709_1), .IN1(~na853_2), .IN2(~na2895_1), .IN3(~na8_2), .IN4(~na3153_1), .IN5(~na2994_1), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y35     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7710_4 ( .OUT(na7710_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7710_6 ( .RAM_O2(na7710_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7710_2), .COMP_OUT(1'b0) );
// C_AND////      x92y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7711_1 ( .OUT(na7711_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7711_6 ( .RAM_O1(na7711_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7711_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7712_4 ( .OUT(na7712_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7712_6 ( .RAM_O2(na7712_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7712_2), .COMP_OUT(1'b0) );
// C_ORAND////      x93y102     80'h00_0018_00_0000_0888_F777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7713_1 ( .OUT(na7713_1), .IN1(~na853_2), .IN2(~na9792_2), .IN3(~na8_2), .IN4(~na3151_1), .IN5(~na9789_2), .IN6(~na1042_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7714_1 ( .OUT(na7714_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7714_6 ( .RAM_O1(na7714_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7714_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7715_4 ( .OUT(na7715_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7715_6 ( .RAM_O2(na7715_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7715_2), .COMP_OUT(1'b0) );
// C_AND////      x92y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7716_1 ( .OUT(na7716_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7716_6 ( .RAM_O1(na7716_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7716_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y48     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7717_4 ( .OUT(na7717_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7717_6 ( .RAM_O2(na7717_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7717_2), .COMP_OUT(1'b0) );
// C_AND////      x92y48     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7718_1 ( .OUT(na7718_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7718_6 ( .RAM_O1(na7718_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7718_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y47     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7719_4 ( .OUT(na7719_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7719_6 ( .RAM_O2(na7719_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7719_2), .COMP_OUT(1'b0) );
// C_AND////      x92y47     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7720_1 ( .OUT(na7720_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7720_6 ( .RAM_O1(na7720_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7720_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y46     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7721_4 ( .OUT(na7721_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7721_6 ( .RAM_O2(na7721_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7721_2), .COMP_OUT(1'b0) );
// C_AND////      x92y46     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7722_1 ( .OUT(na7722_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7722_6 ( .RAM_O1(na7722_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7722_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x77y58     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7723_1 ( .OUT(na7723_1), .IN1(1'b1), .IN2(na9167_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6383_1), .IN8(na6384_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y45     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7724_4 ( .OUT(na7724_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7724_6 ( .RAM_O2(na7724_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7724_2), .COMP_OUT(1'b0) );
// C_AND////      x92y45     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7725_1 ( .OUT(na7725_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7725_6 ( .RAM_O1(na7725_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7725_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y44     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7726_4 ( .OUT(na7726_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7726_6 ( .RAM_O2(na7726_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7726_2), .COMP_OUT(1'b0) );
// C_OR////      x107y68     80'h00_0018_00_0000_0EEE_0DEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7727_1 ( .OUT(na7727_1), .IN1(1'b0), .IN2(na1774_2), .IN3(na1861_2), .IN4(na1464_2), .IN5(~na7728_1), .IN6(na1774_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y67     80'h00_0018_00_0000_0888_4313
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7728_1 ( .OUT(na7728_1), .IN1(1'b1), .IN2(~na1053_2), .IN3(~na1681_1), .IN4(~na7729_2), .IN5(1'b1), .IN6(~na1053_1), .IN7(~na1681_2),
                      .IN8(na1927_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x112y62     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7729_4 ( .OUT(na7729_2), .IN1(na2835_1), .IN2(1'b1), .IN3(na6457_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x109y54     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7730_1 ( .OUT(na7730_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na2942_1), .IN8(~na1921_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7731_1 ( .OUT(na7731_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7731_6 ( .RAM_O1(na7731_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7731_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x89y36     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7732_1 ( .OUT(na7732_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6945_2), .IN8(na7410_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y55     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7733_1 ( .OUT(na7733_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8202_2), .IN8(~na1931_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y43     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7734_4 ( .OUT(na7734_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7734_6 ( .RAM_O2(na7734_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7734_2), .COMP_OUT(1'b0) );
// C_OR////      x105y66     80'h00_0018_00_0000_0EEE_C3EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7735_1 ( .OUT(na7735_1), .IN1(na9533_2), .IN2(1'b0), .IN3(na3140_1), .IN4(na1460_2), .IN5(1'b0), .IN6(~na7736_1), .IN7(1'b0),
                      .IN8(na1770_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y82     80'h00_0018_00_0000_0888_4351
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7736_1 ( .OUT(na7736_1), .IN1(~na7737_2), .IN2(~na1679_1), .IN3(~na1057_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na1679_2), .IN7(~na1057_1),
                      .IN8(na1937_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x111y61     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7737_4 ( .OUT(na7737_2), .IN1(na2835_1), .IN2(1'b1), .IN3(na6458_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x107y54     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7738_1 ( .OUT(na7738_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2941_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1921_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y43     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7739_1 ( .OUT(na7739_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7739_6 ( .RAM_O1(na7739_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7739_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x90y36     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7740_1 ( .OUT(na7740_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7408_1), .IN8(na6944_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y56     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7741_1 ( .OUT(na7741_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1941_1), .IN8(na8201_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7742_4 ( .OUT(na7742_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7742_6 ( .RAM_O2(na7742_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7742_2), .COMP_OUT(1'b0) );
// C_///OR/      x112y52     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7743_4 ( .OUT(na7743_2), .IN1(1'b0), .IN2(~na573_1), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7744_1 ( .OUT(na7744_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7744_6 ( .RAM_O1(na7744_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7744_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x76y56     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7745_1 ( .OUT(na7745_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7451_1), .IN8(na6943_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x100y72     80'h00_0018_00_0000_0EEE_DACA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7746_1 ( .OUT(na7746_1), .IN1(na1607_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1560_2), .IN5(na1607_1), .IN6(1'b0), .IN7(~na7747_1),
                      .IN8(na1579_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y67     80'h00_0018_00_0000_0888_1511
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7747_1 ( .OUT(na7747_1), .IN1(~na1458_1), .IN2(~na1848_2), .IN3(~na1059_2), .IN4(~na1766_2), .IN5(~na1677_2), .IN6(1'b1),
                      .IN7(~na1059_1), .IN8(~na7748_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y62     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7748_1 ( .OUT(na7748_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2835_1), .IN6(1'b1), .IN7(na6461_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y56     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7749_1 ( .OUT(na7749_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1950_1), .IN8(na8200_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7750_4 ( .OUT(na7750_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7750_6 ( .RAM_O2(na7750_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7750_2), .COMP_OUT(1'b0) );
// C_///OR/      x117y50     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7751_4 ( .OUT(na7751_2), .IN1(~na2940_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7752_1 ( .OUT(na7752_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7752_6 ( .RAM_O1(na7752_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7752_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x78y56     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7753_1 ( .OUT(na7753_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6941_1), .IN8(na9957_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x100y66     80'h00_0018_00_0000_0EEE_A3EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7754_1 ( .OUT(na7754_1), .IN1(na1577_2), .IN2(1'b0), .IN3(na1606_2), .IN4(na1558_2), .IN5(1'b0), .IN6(~na7755_1), .IN7(na1606_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y70     80'h00_0018_00_0000_0888_F111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7755_1 ( .OUT(na7755_1), .IN1(~na1846_2), .IN2(~na1747_2), .IN3(~na1443_2), .IN4(~na1761_1), .IN5(~na7756_1), .IN6(~na1747_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y61     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7756_1 ( .OUT(na7756_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2835_1), .IN6(1'b1), .IN7(1'b1), .IN8(na6462_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y54     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7757_1 ( .OUT(na7757_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8736_1), .IN8(~na1959_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7758_1 ( .OUT(na7758_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7758_6 ( .RAM_O1(na7758_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7758_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x115y52     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7759_4 ( .OUT(na7759_2), .IN1(~na2939_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7760_1 ( .OUT(na7760_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7760_6 ( .RAM_O1(na7760_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7760_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x83y86     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7761_1 ( .OUT(na7761_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6984_1), .IN8(na7448_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x85y63     80'h00_0018_00_0000_0EEE_A5EA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7762_1 ( .OUT(na7762_1), .IN1(na1556_2), .IN2(1'b0), .IN3(na1605_2), .IN4(na1575_1), .IN5(~na7763_1), .IN6(1'b0), .IN7(na1605_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x111y71     80'h00_0018_00_0000_0888_F111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7763_1 ( .OUT(na7763_1), .IN1(~na1745_2), .IN2(~na1764_2), .IN3(~na1441_1), .IN4(~na7764_1), .IN5(~na1745_1), .IN6(~na1844_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y64     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7764_1 ( .OUT(na7764_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2835_1), .IN6(1'b1), .IN7(na6465_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y54     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7765_1 ( .OUT(na7765_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8735_2), .IN8(~na1968_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7766_4 ( .OUT(na7766_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7766_6 ( .RAM_O2(na7766_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7766_2), .COMP_OUT(1'b0) );
// C_///OR/      x116y52     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7767_4 ( .OUT(na7767_2), .IN1(~na571_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7768_1 ( .OUT(na7768_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7768_6 ( .RAM_O1(na7768_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7768_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x83y81     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7769_1 ( .OUT(na7769_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6983_2), .IN8(na7447_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x100y71     80'h00_0018_00_0000_0EEE_BCAC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7770_1 ( .OUT(na7770_1), .IN1(1'b0), .IN2(na1599_2), .IN3(na1573_1), .IN4(1'b0), .IN5(1'b0), .IN6(na1599_1), .IN7(na1550_2),
                      .IN8(~na7771_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y74     80'h00_0018_00_0000_0888_F111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7771_1 ( .OUT(na7771_1), .IN1(~na1768_1), .IN2(~na1743_2), .IN3(~na7772_1), .IN4(~na1438_1), .IN5(~na1842_2), .IN6(~na1743_1),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y65     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7772_1 ( .OUT(na7772_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2835_1), .IN6(1'b1), .IN7(na83_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y53     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7773_1 ( .OUT(na7773_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1977_1), .IN8(na8734_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x82y74     80'h00_0078_00_0000_0C88_3AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7774_1 ( .OUT(na7774_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9541_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1984_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7774_4 ( .OUT(na7774_2), .IN1(na7776_1), .IN2(1'b1), .IN3(na977_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y53     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7775_1 ( .OUT(na7775_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1982_1), .IN8(na8733_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y83     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7776_1 ( .OUT(na7776_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7446_1), .IN8(na6982_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7777_4 ( .OUT(na7777_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7777_6 ( .RAM_O2(na7777_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7777_2), .COMP_OUT(1'b0) );
// C_///OR/      x117y48     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7778_4 ( .OUT(na7778_2), .IN1(~na168_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7779_1 ( .OUT(na7779_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7779_6 ( .RAM_O1(na7779_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7779_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x83y69     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7780_1 ( .OUT(na7780_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9541_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1991_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y54     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7781_1 ( .OUT(na7781_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7496_1), .IN8(na6981_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y54     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7782_1 ( .OUT(na7782_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8732_1), .IN8(na1993_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7783_1 ( .OUT(na7783_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7783_6 ( .RAM_O1(na7783_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7783_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x116y50     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7784_4 ( .OUT(na7784_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na170_1), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y43     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7785_1 ( .OUT(na7785_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7785_6 ( .RAM_O1(na7785_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7785_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x102y56     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7786_1 ( .OUT(na7786_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1998_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y56     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7787_1 ( .OUT(na7787_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na6979_1), .IN8(na9958_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y54     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7788_1 ( .OUT(na7788_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8731_2), .IN8(na2000_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7789_4 ( .OUT(na7789_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7789_6 ( .RAM_O2(na7789_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7789_2), .COMP_OUT(1'b0) );
// C_OR////      x110y51     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7790_1 ( .OUT(na7790_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na235_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na1921_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7791_1 ( .OUT(na7791_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7791_6 ( .RAM_O1(na7791_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7791_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x103y54     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7792_1 ( .OUT(na7792_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9541_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na2005_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x55y60     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7793_1 ( .OUT(na7793_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7222_1), .IN8(na7494_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y61     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7794_1 ( .OUT(na7794_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2007_1), .IN8(na8730_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7795_4 ( .OUT(na7795_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7795_6 ( .RAM_O2(na7795_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7795_2), .COMP_OUT(1'b0) );
// C_///OR/      x110y51     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7796_4 ( .OUT(na7796_2), .IN1(1'b0), .IN2(~na246_1), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7797_1 ( .OUT(na7797_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7797_6 ( .RAM_O1(na7797_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7797_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x104y56     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7798_1 ( .OUT(na7798_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9541_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na2012_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y60     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7799_1 ( .OUT(na7799_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7221_2), .IN8(na7484_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y53     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7800_1 ( .OUT(na7800_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2014_1), .IN8(na8729_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x94y48     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7801_4 ( .OUT(na7801_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7801_5 ( .OUT(na7801_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7801_6 ( .RAM_O2(na7801_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7801_2_i), .COMP_OUT(1'b0) );
// C_///OR/      x90y66     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7802_4 ( .OUT(na7802_2), .IN1(~na266_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x94y48     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7803_1 ( .OUT(na7803_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7803_2 ( .OUT(na7803_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7803_6 ( .RAM_O1(na7803_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7803_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x85y71     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7804_1 ( .OUT(na7804_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2019_2), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x56y62     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7805_1 ( .OUT(na7805_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7483_1), .IN8(na7219_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y54     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7806_1 ( .OUT(na7806_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8728_1), .IN8(na2021_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x94y47     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7807_4 ( .OUT(na7807_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7807_5 ( .OUT(na7807_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7807_6 ( .RAM_O2(na7807_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7807_2_i), .COMP_OUT(1'b0) );
// C_///OR/      x107y53     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7808_4 ( .OUT(na7808_2), .IN1(~na269_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x94y47     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7809_1 ( .OUT(na7809_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7809_2 ( .OUT(na7809_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7809_6 ( .RAM_O1(na7809_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7809_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x110y60     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7810_1 ( .OUT(na7810_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9541_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na2026_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y57     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7811_1 ( .OUT(na7811_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7534_1), .IN8(na7218_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y53     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7812_1 ( .OUT(na7812_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8727_2), .IN8(na2028_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y48     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7813_4 ( .OUT(na7813_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7813_5 ( .OUT(na7813_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7813_6 ( .RAM_O2(na7813_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7813_2_i), .COMP_OUT(1'b0) );
// C_///OR/      x109y54     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7814_4 ( .OUT(na7814_2), .IN1(~na270_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y48     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7815_1 ( .OUT(na7815_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7815_2 ( .OUT(na7815_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7815_6 ( .RAM_O1(na7815_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7815_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x106y56     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7816_4 ( .OUT(na7816_2), .IN1(na9541_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2033_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y55     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7817_1 ( .OUT(na7817_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7217_1), .IN8(na9959_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y56     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7818_1 ( .OUT(na7818_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2035_1), .IN8(na8726_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y47     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7819_4 ( .OUT(na7819_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7819_5 ( .OUT(na7819_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7819_6 ( .RAM_O2(na7819_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7819_2_i), .COMP_OUT(1'b0) );
// C_///OR/      x90y62     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7820_4 ( .OUT(na7820_2), .IN1(1'b0), .IN2(~na271_1), .IN3(1'b0), .IN4(~na1921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y47     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7821_1 ( .OUT(na7821_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7821_2 ( .OUT(na7821_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7821_6 ( .RAM_O1(na7821_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7821_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x106y54     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7822_1 ( .OUT(na7822_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2040_1), .IN8(na1921_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y51     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7823_1 ( .OUT(na7823_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7261_1), .IN8(na7531_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y55     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7824_1 ( .OUT(na7824_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2042_1), .IN8(na8725_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y55     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7825_1 ( .OUT(na7825_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8724_1), .IN8(~na2047_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x110y72     80'h00_0060_00_0000_0C0E_FFEA
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7826_4 ( .OUT(na7826_2), .IN1(na1647_2), .IN2(1'b0), .IN3(na1826_2), .IN4(na1722_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y46     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7827_4 ( .OUT(na7827_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7827_5 ( .OUT(na7827_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7827_6 ( .RAM_O2(na7827_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7827_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x108y52     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7828_1 ( .OUT(na7828_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7259_2), .IN8(na7530_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y55     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7829_1 ( .OUT(na7829_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8723_2), .IN8(~na2054_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x106y72     80'h00_0060_00_0000_0C0E_FFEC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7830_4 ( .OUT(na7830_2), .IN1(1'b0), .IN2(na1824_2), .IN3(na1645_2), .IN4(na1720_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y46     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7831_1 ( .OUT(na7831_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7831_2 ( .OUT(na7831_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7831_6 ( .RAM_O1(na7831_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7831_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x107y51     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7832_1 ( .OUT(na7832_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7528_1), .IN8(na7258_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y52     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7833_1 ( .OUT(na7833_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2061_1), .IN8(na8722_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x101y76     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7834_1 ( .OUT(na7834_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1643_1), .IN7(na1822_2), .IN8(na1718_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y45     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7835_4 ( .OUT(na7835_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7835_5 ( .OUT(na7835_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7835_6 ( .RAM_O2(na7835_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7835_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x109y63     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7836_1 ( .OUT(na7836_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7067_1), .IN8(na7257_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y52     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7837_1 ( .OUT(na7837_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2068_1), .IN8(na8721_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x107y72     80'h00_0060_00_0000_0C0E_FFAE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7838_4 ( .OUT(na7838_2), .IN1(na1641_2), .IN2(na1716_2), .IN3(na1820_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y45     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7839_1 ( .OUT(na7839_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7839_2 ( .OUT(na7839_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7839_6 ( .RAM_O1(na7839_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7839_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x110y63     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7840_1 ( .OUT(na7840_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7256_1), .IN8(na9951_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y52     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7841_1 ( .OUT(na7841_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8720_1), .IN8(~na2075_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x108y73     80'h00_0018_00_0000_0CEE_EA00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7842_1 ( .OUT(na7842_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1714_2), .IN6(1'b0), .IN7(na1818_1), .IN8(na1639_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y44     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7843_4 ( .OUT(na7843_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7843_5 ( .OUT(na7843_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7843_6 ( .RAM_O2(na7843_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7843_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x103y63     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7844_1 ( .OUT(na7844_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7329_1), .IN8(na7065_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y52     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7845_1 ( .OUT(na7845_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8719_2), .IN8(~na2082_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y67     80'h00_0018_00_0000_0CEE_AE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7846_1 ( .OUT(na7846_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1712_1), .IN6(na1637_1), .IN7(na1816_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y44     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7847_1 ( .OUT(na7847_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7847_2 ( .OUT(na7847_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7847_6 ( .RAM_O1(na7847_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7847_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x109y62     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7848_1 ( .OUT(na7848_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7328_2), .IN8(na7064_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y55     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7849_1 ( .OUT(na7849_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2089_1), .IN8(na8718_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x103y73     80'h00_0060_00_0000_0C0E_FFAE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7850_4 ( .OUT(na7850_2), .IN1(na1710_2), .IN2(na886_1), .IN3(na1635_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y43     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7851_4 ( .OUT(na7851_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7851_5 ( .OUT(na7851_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7851_6 ( .RAM_O2(na7851_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7851_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x110y62     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7852_1 ( .OUT(na7852_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7061_1), .IN8(na7316_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y51     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7853_1 ( .OUT(na7853_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2096_1), .IN8(na8717_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x103y68     80'h00_0018_00_0000_0CEE_EA00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7854_1 ( .OUT(na7854_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1708_1), .IN6(1'b0), .IN7(na888_2), .IN8(na1633_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y43     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7855_1 ( .OUT(na7855_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7855_2 ( .OUT(na7855_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7855_6 ( .RAM_O1(na7855_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7855_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x100y63     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7856_1 ( .OUT(na7856_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7113_1), .IN8(na7315_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y35     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7857_1 ( .OUT(na7857_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8520_1), .IN8(~na2103_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x105y67     80'h00_0060_00_0000_0C0E_FFCE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7858_4 ( .OUT(na7858_2), .IN1(na1631_1), .IN2(na1706_2), .IN3(1'b0), .IN4(na1814_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y42     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7859_4 ( .OUT(na7859_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7859_5 ( .OUT(na7859_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7859_6 ( .RAM_O2(na7859_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7859_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x103y65     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7860_1 ( .OUT(na7860_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7314_1), .IN8(na9952_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x62y38     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7861_1 ( .OUT(na7861_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8519_2), .IN8(~na2110_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x103y69     80'h00_0060_00_0000_0C0E_FFEC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7862_4 ( .OUT(na7862_2), .IN1(1'b0), .IN2(na1629_2), .IN3(na1704_2), .IN4(na1812_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y42     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7863_1 ( .OUT(na7863_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7863_2 ( .OUT(na7863_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7863_6 ( .RAM_O1(na7863_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7863_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x103y59     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7864_1 ( .OUT(na7864_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7377_1), .IN8(na7110_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x61y40     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7865_1 ( .OUT(na7865_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2117_1), .IN8(na8518_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x104y75     80'h00_0018_00_0000_0CEE_AE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7866_1 ( .OUT(na7866_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1627_1), .IN6(na1702_2), .IN7(na1810_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y41     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7867_4 ( .OUT(na7867_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7867_5 ( .OUT(na7867_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7867_6 ( .RAM_O2(na7867_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7867_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x99y60     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7868_1 ( .OUT(na7868_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7375_2), .IN8(na7107_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x61y38     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7869_1 ( .OUT(na7869_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2124_1), .IN8(na8517_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x99y76     80'h00_0060_00_0000_0C0E_FFEA
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7870_4 ( .OUT(na7870_2), .IN1(na1700_1), .IN2(1'b0), .IN3(na1624_1), .IN4(na1808_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y41     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7871_1 ( .OUT(na7871_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7871_2 ( .OUT(na7871_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7871_6 ( .RAM_O1(na7871_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7871_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x100y62     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7872_1 ( .OUT(na7872_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7105_1), .IN8(na7374_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y58     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7873_1 ( .OUT(na7873_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8516_1), .IN8(~na2131_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x103y68     80'h00_0060_00_0000_0C0E_FFEC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7874_4 ( .OUT(na7874_2), .IN1(1'b0), .IN2(na1698_2), .IN3(na1806_2), .IN4(na1415_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x94y40     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7875_4 ( .OUT(na7875_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7875_5 ( .OUT(na7875_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7875_6 ( .RAM_O2(na7875_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7875_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x81y48     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7876_1 ( .OUT(na7876_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7167_1), .IN8(na7373_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y52     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7877_1 ( .OUT(na7877_1), .IN1(1'b1), .IN2(~na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na8515_2), .IN8(~na2138_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x103y69     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7878_1 ( .OUT(na7878_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1621_2), .IN7(na1691_1), .IN8(na1804_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x94y40     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7879_1 ( .OUT(na7879_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7879_2 ( .OUT(na7879_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7879_6 ( .RAM_O1(na7879_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7879_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x83y49     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7880_1 ( .OUT(na7880_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7370_1), .IN8(na9953_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y40     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7881_1 ( .OUT(na7881_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2145_1), .IN8(na8514_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x104y69     80'h00_0060_00_0000_0C0E_FFCE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7882_4 ( .OUT(na7882_2), .IN1(na1412_2), .IN2(na909_1), .IN3(1'b0), .IN4(na1618_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x94y39     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7883_4 ( .OUT(na7883_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7883_5 ( .OUT(na7883_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7883_6 ( .RAM_O2(na7883_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7883_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x73y43     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7884_1 ( .OUT(na7884_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7414_1), .IN8(na7164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y37     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7885_1 ( .OUT(na7885_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2152_1), .IN8(na8513_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x99y69     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7886_1 ( .OUT(na7886_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1616_1), .IN7(na1689_2), .IN8(na1801_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x94y39     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7887_1 ( .OUT(na7887_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7887_2 ( .OUT(na7887_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7887_6 ( .RAM_O1(na7887_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7887_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x74y44     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7888_1 ( .OUT(na7888_1), .IN1(1'b1), .IN2(na91_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na7412_2), .IN8(na7163_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x128y56     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7889_1 ( .OUT(na7889_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2718_2), .IN7(~na2250_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x57y54     80'h00_0060_00_0000_0C08_FFC4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7890_4 ( .OUT(na7890_2), .IN1(~na3329_2), .IN2(na3263_1), .IN3(1'b1), .IN4(na5961_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x54y46     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7891_4 ( .OUT(na7891_2), .IN1(na3329_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9933_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y40     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7892_4 ( .OUT(na7892_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7892_5 ( .OUT(na7892_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7892_6 ( .RAM_O2(na7892_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7892_2_i), .COMP_OUT(1'b0) );
// C_XOR////      x49y66     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7893_1 ( .OUT(na7893_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na692_1), .IN8(na2311_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y40     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7894_1 ( .OUT(na7894_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7894_2 ( .OUT(na7894_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7894_6 ( .RAM_O1(na7894_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7894_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x49y60     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7895_1 ( .OUT(na7895_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6334_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y39     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7896_4 ( .OUT(na7896_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7896_5 ( .OUT(na7896_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7896_6 ( .RAM_O2(na7896_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7896_2_i), .COMP_OUT(1'b0) );
// C_OR////      x47y58     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7897_1 ( .OUT(na7897_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6333_1), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y39     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7898_1 ( .OUT(na7898_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7898_2 ( .OUT(na7898_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7898_6 ( .RAM_O1(na7898_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7898_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x50y55     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7899_4 ( .OUT(na7899_2), .IN1(~na6327_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y38     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7900_4 ( .OUT(na7900_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7900_5 ( .OUT(na7900_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7900_6 ( .RAM_O2(na7900_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7900_2_i), .COMP_OUT(1'b0) );
// C_OR////      x49y62     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7901_1 ( .OUT(na7901_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6328_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y38     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7902_1 ( .OUT(na7902_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7902_2 ( .OUT(na7902_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7902_6 ( .RAM_O1(na7902_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7902_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x47y54     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7903_1 ( .OUT(na7903_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6317_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y37     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7904_4 ( .OUT(na7904_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7904_5 ( .OUT(na7904_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7904_6 ( .RAM_O2(na7904_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7904_2_i), .COMP_OUT(1'b0) );
// C_///OR/      x49y60     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7905_4 ( .OUT(na7905_2), .IN1(~na6313_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y37     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7906_1 ( .OUT(na7906_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7906_2 ( .OUT(na7906_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7906_6 ( .RAM_O1(na7906_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7906_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y36     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7907_4 ( .OUT(na7907_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7907_5 ( .OUT(na7907_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7907_6 ( .RAM_O2(na7907_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7907_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y36     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7908_1 ( .OUT(na7908_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7908_2 ( .OUT(na7908_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7908_6 ( .RAM_O1(na7908_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7908_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y35     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7909_4 ( .OUT(na7909_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7909_5 ( .OUT(na7909_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7909_6 ( .RAM_O2(na7909_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7909_2_i), .COMP_OUT(1'b0) );
// C_OR////      x47y64     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7910_1 ( .OUT(na7910_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6332_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x96y35     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7911_1 ( .OUT(na7911_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7911_2 ( .OUT(na7911_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7911_6 ( .RAM_O1(na7911_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7911_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR///OR/      x51y55     80'h00_0078_00_0000_0CEE_5757
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7912_1 ( .OUT(na7912_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6325_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7912_4 ( .OUT(na7912_2), .IN1(~na6325_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y34     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7913_4 ( .OUT(na7913_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7913_5 ( .OUT(na7913_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7913_6 ( .RAM_O2(na7913_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7913_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y34     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7914_1 ( .OUT(na7914_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7914_2 ( .OUT(na7914_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7914_6 ( .RAM_O1(na7914_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7914_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y33     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7915_4 ( .OUT(na7915_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7915_5 ( .OUT(na7915_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7915_6 ( .RAM_O2(na7915_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7915_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y33     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7916_1 ( .OUT(na7916_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a7916_2 ( .OUT(na7916_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6645_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7916_6 ( .RAM_O1(na7916_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7916_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y48     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7917_4 ( .OUT(na7917_2), .IN1(1'b1), .IN2(na2878_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7917_6 ( .RAM_O2(na7917_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7917_2), .COMP_OUT(1'b0) );
// C_///OR/      x49y59     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7918_4 ( .OUT(na7918_2), .IN1(~na6315_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y48     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7919_1 ( .OUT(na7919_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2878_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7919_6 ( .RAM_O1(na7919_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7919_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y47     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7920_4 ( .OUT(na7920_2), .IN1(1'b1), .IN2(na2878_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7920_6 ( .RAM_O2(na7920_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7920_2), .COMP_OUT(1'b0) );
// C_AND////      x93y47     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7921_1 ( .OUT(na7921_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2878_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7921_6 ( .RAM_O1(na7921_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7921_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x50y55     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7922_1 ( .OUT(na7922_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9806_2), .IN6(~na369_2), .IN7(~na6314_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y48     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7923_4 ( .OUT(na7923_2), .IN1(1'b1), .IN2(na2878_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7923_6 ( .RAM_O2(na7923_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7923_2), .COMP_OUT(1'b0) );
// C_///OR/      x52y57     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7924_4 ( .OUT(na7924_2), .IN1(~na6331_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y48     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7925_1 ( .OUT(na7925_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2878_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7925_6 ( .RAM_O1(na7925_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7925_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR///OR/      x49y57     80'h00_0078_00_0000_0CEE_5757
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7926_1 ( .OUT(na7926_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6320_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7926_4 ( .OUT(na7926_2), .IN1(~na6320_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y47     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7927_4 ( .OUT(na7927_2), .IN1(1'b1), .IN2(na2878_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7927_6 ( .RAM_O2(na7927_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7927_2), .COMP_OUT(1'b0) );
// C_OR////      x49y59     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7928_1 ( .OUT(na7928_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na9806_2), .IN6(~na369_2), .IN7(~na6330_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y47     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7929_1 ( .OUT(na7929_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2878_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7929_6 ( .RAM_O1(na7929_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7929_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x57y63     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7930_4 ( .OUT(na7930_2), .IN1(~na6336_2), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y46     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7931_4 ( .OUT(na7931_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2877_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7931_6 ( .RAM_O2(na7931_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7931_2), .COMP_OUT(1'b0) );
// C_AND////      x95y46     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7932_1 ( .OUT(na7932_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2877_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7932_6 ( .RAM_O1(na7932_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7932_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y45     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7933_4 ( .OUT(na7933_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2877_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7933_6 ( .RAM_O2(na7933_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7933_2), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x48y62     80'h00_0078_00_0000_0C66_60AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7934_1 ( .OUT(na7934_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2357_2), .IN8(na612_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7934_4 ( .OUT(na7934_2), .IN1(na1586_1), .IN2(1'b0), .IN3(na2357_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y45     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7935_1 ( .OUT(na7935_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2877_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7935_6 ( .RAM_O1(na7935_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7935_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x49y53     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7936_1 ( .OUT(na7936_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6326_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y44     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7937_4 ( .OUT(na7937_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2877_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7937_6 ( .RAM_O2(na7937_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7937_2), .COMP_OUT(1'b0) );
// C_///OR/      x47y54     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7938_4 ( .OUT(na7938_2), .IN1(~na6319_2), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y44     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7939_1 ( .OUT(na7939_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2877_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7939_6 ( .RAM_O1(na7939_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7939_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x49y53     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7940_4 ( .OUT(na7940_2), .IN1(~na6312_2), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y43     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7941_4 ( .OUT(na7941_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2877_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7941_6 ( .RAM_O2(na7941_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7941_2), .COMP_OUT(1'b0) );
// C_///OR/      x49y58     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7942_4 ( .OUT(na7942_2), .IN1(~na9806_2), .IN2(~na369_2), .IN3(~na6329_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y43     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7943_1 ( .OUT(na7943_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2877_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7943_6 ( .RAM_O1(na7943_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7943_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x48y60     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7944_1 ( .OUT(na7944_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6323_1), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y42     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7945_4 ( .OUT(na7945_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2876_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7945_6 ( .RAM_O2(na7945_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7945_2), .COMP_OUT(1'b0) );
// C_AND////      x95y42     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7946_1 ( .OUT(na7946_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2876_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7946_6 ( .RAM_O1(na7946_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7946_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y41     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7947_4 ( .OUT(na7947_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2876_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7947_6 ( .RAM_O2(na7947_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7947_2), .COMP_OUT(1'b0) );
// C_OR///OR/      x50y53     80'h00_0078_00_0000_0CEE_5757
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7948_1 ( .OUT(na7948_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6324_2), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7948_4 ( .OUT(na7948_2), .IN1(~na6324_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y41     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7949_1 ( .OUT(na7949_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2876_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7949_6 ( .RAM_O1(na7949_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7949_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x48y58     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7950_4 ( .OUT(na7950_2), .IN1(~na6318_1), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y40     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7951_4 ( .OUT(na7951_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2853_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7951_6 ( .RAM_O2(na7951_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7951_2), .COMP_OUT(1'b0) );
// C_///XOR/      x50y63     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7952_4 ( .OUT(na7952_2), .IN1(na2383_2), .IN2(1'b0), .IN3(1'b0), .IN4(na617_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x47y62     80'h00_0078_00_0000_0C66_CAAA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7953_1 ( .OUT(na7953_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na50_2), .IN6(1'b0), .IN7(1'b0), .IN8(na355_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7953_4 ( .OUT(na7953_2), .IN1(na2383_1), .IN2(1'b0), .IN3(na627_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x50y64     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7954_1 ( .OUT(na7954_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na50_1), .IN6(1'b0), .IN7(na357_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x51y67     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7955_1 ( .OUT(na7955_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2385_1), .IN6(1'b0), .IN7(1'b0), .IN8(na702_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y40     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7956_1 ( .OUT(na7956_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2853_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7956_6 ( .RAM_O1(na7956_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7956_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x50y52     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a7957_4 ( .OUT(na7957_2), .IN1(~na6322_2), .IN2(~na369_2), .IN3(~na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y39     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7958_4 ( .OUT(na7958_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2853_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7958_6 ( .RAM_O2(na7958_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7958_2), .COMP_OUT(1'b0) );
// C_OR////      x49y58     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7959_1 ( .OUT(na7959_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6335_1), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y39     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7960_1 ( .OUT(na7960_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2853_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7960_6 ( .RAM_O1(na7960_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7960_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x45y52     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a7961_1 ( .OUT(na7961_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na6321_1), .IN6(~na369_2), .IN7(~na3268_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y40     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7962_4 ( .OUT(na7962_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2853_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7962_6 ( .RAM_O2(na7962_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7962_2), .COMP_OUT(1'b0) );
// C_ORAND////      x84y59     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7963_1 ( .OUT(na7963_1), .IN1(na7966_2), .IN2(na9545_2), .IN3(~na10016_2), .IN4(1'b0), .IN5(~na7966_2), .IN6(na9555_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y40     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7964_1 ( .OUT(na7964_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2853_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7964_6 ( .RAM_O1(na7964_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7964_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y39     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7965_4 ( .OUT(na7965_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2853_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7965_6 ( .RAM_O2(na7965_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7965_2), .COMP_OUT(1'b0) );
// C_AND///AND/      x85y37     80'h00_0078_00_0000_0C88_555A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7966_1 ( .OUT(na7966_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na5692_2), .IN6(1'b1), .IN7(~na5691_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7966_4 ( .OUT(na7966_2), .IN1(na5692_1), .IN2(1'b1), .IN3(~na5691_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y39     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7967_1 ( .OUT(na7967_1), .IN1(na7966_2), .IN2(na9546_2), .IN3(~na10016_2), .IN4(1'b0), .IN5(~na7966_2), .IN6(na9556_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y39     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7968_1 ( .OUT(na7968_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2853_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7968_6 ( .RAM_O1(na7968_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7968_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y38     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7969_4 ( .OUT(na7969_2), .IN1(na2850_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7969_6 ( .RAM_O2(na7969_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7969_2), .COMP_OUT(1'b0) );
// C_AND////      x95y38     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7970_1 ( .OUT(na7970_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2850_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7970_6 ( .RAM_O1(na7970_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7970_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x86y40     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7971_1 ( .OUT(na7971_1), .IN1(na7966_2), .IN2(na9547_2), .IN3(~na10016_2), .IN4(1'b0), .IN5(~na7966_2), .IN6(na9557_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y37     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7972_4 ( .OUT(na7972_2), .IN1(na2850_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7972_6 ( .RAM_O2(na7972_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7972_2), .COMP_OUT(1'b0) );
// C_AND////      x95y37     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7973_1 ( .OUT(na7973_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2850_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7973_6 ( .RAM_O1(na7973_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7973_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y36     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7974_4 ( .OUT(na7974_2), .IN1(na2850_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7974_6 ( .RAM_O2(na7974_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7974_2), .COMP_OUT(1'b0) );
// C_ORAND////      x83y40     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7975_1 ( .OUT(na7975_1), .IN1(na7966_2), .IN2(na2008_2), .IN3(~na10016_2), .IN4(1'b0), .IN5(~na7966_2), .IN6(na9558_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y36     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7976_1 ( .OUT(na7976_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2850_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7976_6 ( .RAM_O1(na7976_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7976_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y35     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7977_4 ( .OUT(na7977_2), .IN1(na2850_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7977_6 ( .RAM_O2(na7977_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7977_2), .COMP_OUT(1'b0) );
// C_AND////      x95y35     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7978_1 ( .OUT(na7978_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2850_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7978_6 ( .RAM_O1(na7978_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7978_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x88y42     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7979_1 ( .OUT(na7979_1), .IN1(na7966_2), .IN2(na9549_2), .IN3(~na10016_2), .IN4(1'b0), .IN5(~na7966_2), .IN6(na9559_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y34     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7980_4 ( .OUT(na7980_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2846_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7980_6 ( .RAM_O2(na7980_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7980_2), .COMP_OUT(1'b0) );
// C_AND////      x95y34     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7981_1 ( .OUT(na7981_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2846_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7981_6 ( .RAM_O1(na7981_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7981_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y33     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7982_4 ( .OUT(na7982_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2846_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7982_6 ( .RAM_O2(na7982_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7982_2), .COMP_OUT(1'b0) );
// C_ORAND////      x86y44     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7983_1 ( .OUT(na7983_1), .IN1(na7966_2), .IN2(na9550_2), .IN3(~na10016_2), .IN4(1'b0), .IN5(~na7966_2), .IN6(na9560_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y33     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7984_1 ( .OUT(na7984_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2846_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7984_6 ( .RAM_O1(na7984_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7984_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x99y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7985_1 ( .OUT(na7985_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7985_6 ( .RAM_O1(na7985_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7985_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x91y65     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7986_4 ( .OUT(na7986_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3242_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7986_6 ( .RAM_O2(na7986_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7986_2), .COMP_OUT(1'b0) );
// C_ORAND////      x88y44     80'h00_0018_00_0000_0888_FD5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7987_1 ( .OUT(na7987_1), .IN1(na7966_2), .IN2(na9551_2), .IN3(~na10016_2), .IN4(1'b0), .IN5(~na7966_2), .IN6(na9562_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y72     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7988_4 ( .OUT(na7988_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7988_6 ( .RAM_O2(na7988_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7988_2), .COMP_OUT(1'b0) );
// C_AND////      x92y72     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7989_1 ( .OUT(na7989_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7989_6 ( .RAM_O1(na7989_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7989_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y71     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7990_4 ( .OUT(na7990_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7990_6 ( .RAM_O2(na7990_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7990_2), .COMP_OUT(1'b0) );
// C_AND////      x92y71     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7991_1 ( .OUT(na7991_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7991_6 ( .RAM_O1(na7991_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7991_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y70     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7992_4 ( .OUT(na7992_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7992_6 ( .RAM_O2(na7992_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7992_2), .COMP_OUT(1'b0) );
// C_AND////      x92y70     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7993_1 ( .OUT(na7993_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7993_6 ( .RAM_O1(na7993_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7993_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x79y63     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7994_4 ( .OUT(na7994_2), .IN1(na5692_2), .IN2(na2043_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y69     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7995_4 ( .OUT(na7995_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7995_6 ( .RAM_O2(na7995_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7995_2), .COMP_OUT(1'b0) );
// C_AND////      x92y69     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7996_1 ( .OUT(na7996_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7996_6 ( .RAM_O1(na7996_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7996_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x73y61     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7997_1 ( .OUT(na7997_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(na2050_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y68     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7998_4 ( .OUT(na7998_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7998_6 ( .RAM_O2(na7998_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na7998_2), .COMP_OUT(1'b0) );
// C_AND////      x92y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7999_1 ( .OUT(na7999_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a7999_6 ( .RAM_O1(na7999_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na7999_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x79y59     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8000_1 ( .OUT(na8000_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(na2057_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y67     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8001_4 ( .OUT(na8001_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8001_6 ( .RAM_O2(na8001_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8001_2), .COMP_OUT(1'b0) );
// C_AND////      x92y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8002_1 ( .OUT(na8002_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8002_6 ( .RAM_O1(na8002_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8002_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x81y59     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8003_1 ( .OUT(na8003_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2064_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8004_4 ( .OUT(na8004_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8004_6 ( .RAM_O2(na8004_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8004_2), .COMP_OUT(1'b0) );
// C_AND////      x92y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8005_1 ( .OUT(na8005_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8005_6 ( .RAM_O1(na8005_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8005_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y57     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8006_4 ( .OUT(na8006_2), .IN1(na5692_2), .IN2(na2071_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8007_4 ( .OUT(na8007_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8007_6 ( .RAM_O2(na8007_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8007_2), .COMP_OUT(1'b0) );
// C_AND////      x92y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8008_1 ( .OUT(na8008_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8008_6 ( .RAM_O1(na8008_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8008_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x83y55     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8009_1 ( .OUT(na8009_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2078_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8010_1 ( .OUT(na8010_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8010_6 ( .RAM_O1(na8010_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8010_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x101y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8011_1 ( .OUT(na8011_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8011_6 ( .RAM_O1(na8011_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8011_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x73y57     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8012_1 ( .OUT(na8012_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(na2085_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8013_4 ( .OUT(na8013_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8013_6 ( .RAM_O2(na8013_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8013_2), .COMP_OUT(1'b0) );
// C_AND////      x101y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8014_1 ( .OUT(na8014_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8014_6 ( .RAM_O1(na8014_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8014_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x75y59     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8015_1 ( .OUT(na8015_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(na2092_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8016_4 ( .OUT(na8016_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8016_6 ( .RAM_O2(na8016_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8016_2), .COMP_OUT(1'b0) );
// C_AND////      x101y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8017_1 ( .OUT(na8017_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8017_6 ( .RAM_O1(na8017_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8017_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x83y43     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8018_4 ( .OUT(na8018_2), .IN1(na5692_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2099_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x94y72     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8019_4 ( .OUT(na8019_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8019_5 ( .OUT(na8019_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8019_6 ( .RAM_O2(na8019_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8019_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x94y72     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8020_1 ( .OUT(na8020_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8020_2 ( .OUT(na8020_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8020_6 ( .RAM_O1(na8020_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8020_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x73y59     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8021_1 ( .OUT(na8021_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2106_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x94y71     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8022_4 ( .OUT(na8022_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8022_5 ( .OUT(na8022_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8022_6 ( .RAM_O2(na8022_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8022_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x94y71     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8023_1 ( .OUT(na8023_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8023_2 ( .OUT(na8023_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8023_6 ( .RAM_O1(na8023_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8023_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x83y45     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8024_4 ( .OUT(na8024_2), .IN1(na5692_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2113_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y72     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8025_4 ( .OUT(na8025_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8025_5 ( .OUT(na8025_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8025_6 ( .RAM_O2(na8025_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8025_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y72     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8026_1 ( .OUT(na8026_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8026_2 ( .OUT(na8026_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8026_6 ( .RAM_O1(na8026_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8026_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x81y49     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8027_1 ( .OUT(na8027_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2120_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y71     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8028_4 ( .OUT(na8028_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8028_5 ( .OUT(na8028_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8028_6 ( .RAM_O2(na8028_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8028_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y71     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8029_1 ( .OUT(na8029_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8029_2 ( .OUT(na8029_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8029_6 ( .RAM_O1(na8029_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8029_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x83y47     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8030_4 ( .OUT(na8030_2), .IN1(na5692_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2127_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y70     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8031_4 ( .OUT(na8031_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8031_5 ( .OUT(na8031_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8031_6 ( .RAM_O2(na8031_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8031_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y70     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8032_1 ( .OUT(na8032_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8032_2 ( .OUT(na8032_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8032_6 ( .RAM_O1(na8032_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8032_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x81y51     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8033_1 ( .OUT(na8033_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2134_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y69     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8034_4 ( .OUT(na8034_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8034_5 ( .OUT(na8034_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8034_6 ( .RAM_O2(na8034_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8034_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y69     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8035_1 ( .OUT(na8035_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8035_2 ( .OUT(na8035_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8035_6 ( .RAM_O1(na8035_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8035_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x81y45     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8036_4 ( .OUT(na8036_2), .IN1(na5692_2), .IN2(1'b1), .IN3(1'b1), .IN4(na2141_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y68     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8037_4 ( .OUT(na8037_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8037_5 ( .OUT(na8037_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8037_6 ( .RAM_O2(na8037_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8037_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y68     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8038_1 ( .OUT(na8038_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8038_2 ( .OUT(na8038_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8038_6 ( .RAM_O1(na8038_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8038_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x81y47     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8039_1 ( .OUT(na8039_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na5692_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2148_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x96y67     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8040_4 ( .OUT(na8040_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8040_5 ( .OUT(na8040_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8040_6 ( .RAM_O2(na8040_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8040_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y67     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8041_1 ( .OUT(na8041_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8041_2 ( .OUT(na8041_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8041_6 ( .RAM_O1(na8041_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8041_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y66     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8042_4 ( .OUT(na8042_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8042_5 ( .OUT(na8042_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8042_6 ( .RAM_O2(na8042_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8042_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y66     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8043_1 ( .OUT(na8043_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8043_2 ( .OUT(na8043_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8043_6 ( .RAM_O1(na8043_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8043_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y65     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8044_4 ( .OUT(na8044_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8044_5 ( .OUT(na8044_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8044_6 ( .RAM_O2(na8044_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8044_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y65     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8045_1 ( .OUT(na8045_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8045_2 ( .OUT(na8045_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6647_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8045_6 ( .RAM_O1(na8045_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8045_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y72     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8046_4 ( .OUT(na8046_2), .IN1(na2885_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8046_6 ( .RAM_O2(na8046_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8046_2), .COMP_OUT(1'b0) );
// C_AND////      x93y72     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8047_1 ( .OUT(na8047_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2885_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8047_6 ( .RAM_O1(na8047_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8047_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y71     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8048_4 ( .OUT(na8048_2), .IN1(na2885_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8048_6 ( .RAM_O2(na8048_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8048_2), .COMP_OUT(1'b0) );
// C_AND////      x93y71     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8049_1 ( .OUT(na8049_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2885_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8049_6 ( .RAM_O1(na8049_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8049_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y72     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8050_4 ( .OUT(na8050_2), .IN1(na2885_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8050_6 ( .RAM_O2(na8050_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8050_2), .COMP_OUT(1'b0) );
// C_AND////      x95y72     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8051_1 ( .OUT(na8051_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2885_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8051_6 ( .RAM_O1(na8051_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8051_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y71     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8052_4 ( .OUT(na8052_2), .IN1(na2885_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8052_6 ( .RAM_O2(na8052_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8052_2), .COMP_OUT(1'b0) );
// C_AND////      x95y71     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8053_1 ( .OUT(na8053_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2885_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8053_6 ( .RAM_O1(na8053_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8053_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y70     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8054_4 ( .OUT(na8054_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8054_6 ( .RAM_O2(na8054_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8054_2), .COMP_OUT(1'b0) );
// C_AND////      x95y70     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8055_1 ( .OUT(na8055_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8055_6 ( .RAM_O1(na8055_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8055_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y69     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8056_4 ( .OUT(na8056_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8056_6 ( .RAM_O2(na8056_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8056_2), .COMP_OUT(1'b0) );
// C_AND////      x95y69     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8057_1 ( .OUT(na8057_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8057_6 ( .RAM_O1(na8057_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8057_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x119y100     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8058_4 ( .OUT(na8058_2), .IN1(1'b1), .IN2(na1064_1), .IN3(na9369_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y68     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8059_4 ( .OUT(na8059_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8059_6 ( .RAM_O2(na8059_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8059_2), .COMP_OUT(1'b0) );
// C_AND////      x95y68     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8060_1 ( .OUT(na8060_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8060_6 ( .RAM_O1(na8060_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8060_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x127y75     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8061_1 ( .OUT(na8061_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2706_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y67     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8062_4 ( .OUT(na8062_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2883_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8062_6 ( .RAM_O2(na8062_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8062_2), .COMP_OUT(1'b0) );
// C_///AND/      x129y66     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8063_4 ( .OUT(na8063_2), .IN1(~na296_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2708_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y67     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8064_1 ( .OUT(na8064_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2883_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8064_6 ( .RAM_O1(na8064_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8064_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x129y68     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8065_4 ( .OUT(na8065_2), .IN1(~na296_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2710_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y66     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8066_4 ( .OUT(na8066_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2882_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8066_6 ( .RAM_O2(na8066_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8066_2), .COMP_OUT(1'b0) );
// C_///AND/      x131y68     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8067_4 ( .OUT(na8067_2), .IN1(~na296_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2712_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y66     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8068_1 ( .OUT(na8068_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2882_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8068_6 ( .RAM_O1(na8068_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8068_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x123y69     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8069_1 ( .OUT(na8069_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2714_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x132y52     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8070_4 ( .OUT(na8070_2), .IN1(na3881_2), .IN2(1'b1), .IN3(~na2250_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y65     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8071_4 ( .OUT(na8071_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2882_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8071_6 ( .RAM_O2(na8071_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8071_2), .COMP_OUT(1'b0) );
// C_AND////      x127y71     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8072_1 ( .OUT(na8072_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2723_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y99     80'h00_0060_00_0000_0C08_FFA2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8073_4 ( .OUT(na8073_2), .IN1(na1039_1), .IN2(~na6065_2), .IN3(na953_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y65     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8074_1 ( .OUT(na8074_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2882_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8074_6 ( .RAM_O1(na8074_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8074_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x127y61     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8075_4 ( .OUT(na8075_2), .IN1(~na296_1), .IN2(1'b1), .IN3(na2735_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x132y52     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8076_1 ( .OUT(na8076_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3881_1), .IN6(1'b1), .IN7(~na2250_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x133y52     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8077_4 ( .OUT(na8077_2), .IN1(1'b1), .IN2(na3883_1), .IN3(~na2250_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y69     80'h00_0018_00_0000_0C88_A4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8078_1 ( .OUT(na8078_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6118_2), .IN6(na2834_1), .IN7(na2808_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y89     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8079_1 ( .OUT(na8079_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8079_6 ( .RAM_O1(na8079_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8079_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x125y75     80'h00_0018_00_0000_0C88_BCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8080_1 ( .OUT(na8080_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na2768_2), .IN7(na2770_1), .IN8(~na8081_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x130y74     80'h00_0060_00_0000_0C0E_FFAE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a8081_4 ( .OUT(na8081_2), .IN1(na6936_2), .IN2(na99_2), .IN3(na298_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8082_1 ( .OUT(na8082_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8082_6 ( .RAM_O1(na8082_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8082_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x59y89     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8083_4 ( .OUT(na8083_2), .IN1(1'b1), .IN2(na3241_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8083_6 ( .RAM_O2(na8083_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8083_2), .COMP_OUT(1'b0) );
// C_///AND/      x59y81     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8084_4 ( .OUT(na8084_2), .IN1(1'b1), .IN2(na3248_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8084_6 ( .RAM_O2(na8084_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8084_2), .COMP_OUT(1'b0) );
// C_MX4b////      x77y82     80'h00_0018_00_0040_0A68_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a8085_1 ( .OUT(na8085_1), .IN1(~na712_1), .IN2(1'b1), .IN3(1'b1), .IN4(na523_1), .IN5(1'b0), .IN6(na2773_1), .IN7(na9674_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y88     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8086_4 ( .OUT(na8086_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8086_6 ( .RAM_O2(na8086_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8086_2), .COMP_OUT(1'b0) );
// C_AND////      x123y72     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8087_1 ( .OUT(na8087_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2774_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y88     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8088_1 ( .OUT(na8088_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8088_6 ( .RAM_O1(na8088_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8088_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x121y72     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8089_1 ( .OUT(na8089_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2776_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y87     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8090_4 ( .OUT(na8090_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8090_6 ( .RAM_O2(na8090_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8090_2), .COMP_OUT(1'b0) );
// C_AND////      x131y74     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8091_1 ( .OUT(na8091_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na296_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2778_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x130y51     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8092_4 ( .OUT(na8092_2), .IN1(~na985_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na989_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x135y96     80'h00_0018_00_0000_0888_F5B3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8093_1 ( .OUT(na8093_1), .IN1(1'b0), .IN2(~na215_1), .IN3(na8094_1), .IN4(~na2836_2), .IN5(~na6936_2), .IN6(1'b0), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x124y91     80'h00_0018_00_0000_0888_A82A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8094_1 ( .OUT(na8094_1), .IN1(na652_1), .IN2(1'b1), .IN3(na709_2), .IN4(~na753_1), .IN5(na652_2), .IN6(na2894_2), .IN7(na2838_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x73y54     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8095_1 ( .OUT(na8095_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na356_2), .IN6(1'b1), .IN7(~na354_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y55     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8096_4 ( .OUT(na8096_2), .IN1(1'b1), .IN2(~na5402_1), .IN3(1'b1), .IN4(~na5403_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x83y50     80'h00_0060_00_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a8097_4 ( .OUT(na8097_2), .IN1(1'b0), .IN2(~na798_2), .IN3(na354_2), .IN4(na5403_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y75     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8098_1 ( .OUT(na8098_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na354_2), .IN8(~na5403_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x127y99     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8099_4 ( .OUT(na8099_2), .IN1(1'b0), .IN2(na2919_1), .IN3(na106_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y87     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8100_1 ( .OUT(na8100_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8100_6 ( .RAM_O1(na8100_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8100_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x136y65     80'h00_0078_00_0000_0C88_C315
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8101_1 ( .OUT(na8101_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na6475_1), .IN7(1'b1), .IN8(na154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8101_4 ( .OUT(na8101_2), .IN1(~na1010_1), .IN2(1'b1), .IN3(~na1016_1), .IN4(~na1018_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y86     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8102_4 ( .OUT(na8102_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8102_6 ( .RAM_O2(na8102_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8102_2), .COMP_OUT(1'b0) );
// C_AND////      x125y91     80'h00_0018_00_0000_0888_5A2A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8103_1 ( .OUT(na8103_1), .IN1(na652_1), .IN2(1'b1), .IN3(na224_1), .IN4(~na753_1), .IN5(na652_2), .IN6(1'b1), .IN7(~na709_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x87y91     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8104_1 ( .OUT(na8104_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2935_1), .IN7(na2937_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y86     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8105_1 ( .OUT(na8105_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8105_6 ( .RAM_O1(na8105_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8105_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x120y52     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8106_1 ( .OUT(na8106_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8107_2), .IN6(1'b1), .IN7(na2950_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x123y53     80'h00_0078_00_0000_0C88_5C35
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8107_1 ( .OUT(na8107_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2921_1), .IN7(~na2950_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8107_4 ( .OUT(na8107_2), .IN1(~na10027_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y85     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8108_4 ( .OUT(na8108_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8108_6 ( .RAM_O2(na8108_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8108_2), .COMP_OUT(1'b0) );
// C_///AND/      x119y97     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8109_4 ( .OUT(na8109_2), .IN1(na2951_2), .IN2(1'b1), .IN3(1'b1), .IN4(na9296_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y85     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8110_1 ( .OUT(na8110_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8110_6 ( .RAM_O1(na8110_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8110_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x123y95     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8111_4 ( .OUT(na8111_2), .IN1(na643_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2953_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y84     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8112_4 ( .OUT(na8112_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8112_6 ( .RAM_O2(na8112_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8112_2), .COMP_OUT(1'b0) );
// C_AND////      x125y93     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8113_1 ( .OUT(na8113_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na643_1), .IN6(1'b1), .IN7(1'b1), .IN8(na753_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y84     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8114_1 ( .OUT(na8114_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8114_6 ( .RAM_O1(na8114_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8114_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y83     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8115_4 ( .OUT(na8115_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8115_6 ( .RAM_O2(na8115_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8115_2), .COMP_OUT(1'b0) );
// C_///AND/      x132y46     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8116_4 ( .OUT(na8116_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3888_2), .IN4(~na989_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y83     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8117_1 ( .OUT(na8117_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8117_6 ( .RAM_O1(na8117_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8117_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x115y63     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8118_1 ( .OUT(na8118_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2981_1), .IN6(~na9186_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x116y102     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8119_4 ( .OUT(na8119_2), .IN1(na2987_1), .IN2(~na2983_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y82     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8120_4 ( .OUT(na8120_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8120_6 ( .RAM_O2(na8120_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8120_2), .COMP_OUT(1'b0) );
// C_OR////      x118y98     80'h00_0018_00_0000_0CEE_D300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8121_1 ( .OUT(na8121_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1064_2), .IN7(~na9387_2), .IN8(na238_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8122_1 ( .OUT(na8122_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8122_6 ( .RAM_O1(na8122_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8122_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR////      x121y100     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8123_1 ( .OUT(na8123_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2987_1), .IN6(1'b0), .IN7(1'b0), .IN8(na2984_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8124_4 ( .OUT(na8124_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8124_6 ( .RAM_O2(na8124_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8124_2), .COMP_OUT(1'b0) );
// C_///AND/      x101y67     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8125_4 ( .OUT(na8125_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1132_1), .IN4(~na2980_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8126_1 ( .OUT(na8126_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8126_6 ( .RAM_O1(na8126_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8126_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y96     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8127_4 ( .OUT(na8127_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8127_6 ( .RAM_O2(na8127_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8127_2), .COMP_OUT(1'b0) );
// C_AND////      x60y96     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8128_1 ( .OUT(na8128_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8128_6 ( .RAM_O1(na8128_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8128_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y95     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8129_4 ( .OUT(na8129_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8129_6 ( .RAM_O2(na8129_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8129_2), .COMP_OUT(1'b0) );
// C_AND////      x107y59     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8130_1 ( .OUT(na8130_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na9412_2), .IN7(1'b1), .IN8(na1135_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y95     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8131_1 ( .OUT(na8131_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8131_6 ( .RAM_O1(na8131_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8131_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x109y59     80'h00_0078_00_0000_0C88_8F8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8132_1 ( .OUT(na8132_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1165_2), .IN8(na1135_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8132_4 ( .OUT(na8132_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1165_1), .IN4(na1135_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y94     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8133_4 ( .OUT(na8133_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8133_6 ( .RAM_O2(na8133_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8133_2), .COMP_OUT(1'b0) );
// C_///AND/      x125y75     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8134_4 ( .OUT(na8134_2), .IN1(1'b1), .IN2(~na3029_2), .IN3(na9510_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y94     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8135_1 ( .OUT(na8135_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8135_6 ( .RAM_O1(na8135_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8135_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y93     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8136_4 ( .OUT(na8136_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8136_6 ( .RAM_O2(na8136_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8136_2), .COMP_OUT(1'b0) );
// C_AND////      x94y99     80'h00_0018_00_0000_0C88_2AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8137_1 ( .OUT(na8137_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3354_1), .IN6(1'b1), .IN7(na3276_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y93     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8138_1 ( .OUT(na8138_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8138_6 ( .RAM_O1(na8138_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8138_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y92     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8139_4 ( .OUT(na8139_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8139_6 ( .RAM_O2(na8139_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8139_2), .COMP_OUT(1'b0) );
// C_AND////      x60y92     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8140_1 ( .OUT(na8140_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8140_6 ( .RAM_O1(na8140_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8140_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y91     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8141_4 ( .OUT(na8141_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8141_6 ( .RAM_O2(na8141_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8141_2), .COMP_OUT(1'b0) );
// C_OR////      x116y72     80'h00_0018_00_0000_0CEE_3B00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8142_1 ( .OUT(na8142_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3225_1), .IN6(~na3222_1), .IN7(1'b0), .IN8(~na3226_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y91     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8143_1 ( .OUT(na8143_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8143_6 ( .RAM_O1(na8143_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8143_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y90     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8144_4 ( .OUT(na8144_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8144_6 ( .RAM_O2(na8144_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8144_2), .COMP_OUT(1'b0) );
// C_AND////      x60y90     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8145_1 ( .OUT(na8145_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8145_6 ( .RAM_O1(na8145_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8145_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y89     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8146_4 ( .OUT(na8146_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8146_6 ( .RAM_O2(na8146_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8146_2), .COMP_OUT(1'b0) );
// C_AND////      x60y89     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8147_1 ( .OUT(na8147_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8147_6 ( .RAM_O1(na8147_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8147_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y84     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8148_1 ( .OUT(na8148_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8148_6 ( .RAM_O1(na8148_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8148_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y83     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8149_1 ( .OUT(na8149_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8149_6 ( .RAM_O1(na8149_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8149_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y82     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8150_4 ( .OUT(na8150_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8150_6 ( .RAM_O2(na8150_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8150_2), .COMP_OUT(1'b0) );
// C_XOR////      x130y118     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8151_1 ( .OUT(na8151_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na6055_1), .IN6(~na318_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x129y116     80'h00_0060_00_0000_0C06_FF5A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8152_4 ( .OUT(na8152_2), .IN1(na6055_1), .IN2(1'b0), .IN3(~na320_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8153_1 ( .OUT(na8153_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8153_6 ( .RAM_O1(na8153_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8153_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x115y103     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8154_1 ( .OUT(na8154_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1039_1), .IN6(1'b1), .IN7(na953_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8155_4 ( .OUT(na8155_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8155_6 ( .RAM_O2(na8155_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8155_2), .COMP_OUT(1'b0) );
// C_AND////      x69y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8156_1 ( .OUT(na8156_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8156_6 ( .RAM_O1(na8156_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8156_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y92     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8157_1 ( .OUT(na8157_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8157_6 ( .RAM_O1(na8157_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8157_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x123y62     80'h00_0018_00_0000_0888_3FEA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8158_1 ( .OUT(na8158_1), .IN1(na3225_1), .IN2(1'b0), .IN3(na9798_2), .IN4(na3227_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(~na6626_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y91     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8159_1 ( .OUT(na8159_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8159_6 ( .RAM_O1(na8159_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8159_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y90     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8160_4 ( .OUT(na8160_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8160_6 ( .RAM_O2(na8160_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8160_2), .COMP_OUT(1'b0) );
// C_AND////      x69y90     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8161_1 ( .OUT(na8161_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8161_6 ( .RAM_O1(na8161_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8161_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y89     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8162_4 ( .OUT(na8162_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8162_6 ( .RAM_O2(na8162_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8162_2), .COMP_OUT(1'b0) );
// C_AND////      x69y89     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8163_1 ( .OUT(na8163_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8163_6 ( .RAM_O1(na8163_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8163_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y96     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8164_4 ( .OUT(na8164_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8164_5 ( .OUT(na8164_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8164_6 ( .RAM_O2(na8164_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8164_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y96     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8165_1 ( .OUT(na8165_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8165_2 ( .OUT(na8165_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8165_6 ( .RAM_O1(na8165_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8165_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x111y68     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8166_1 ( .OUT(na8166_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2834_1), .IN7(na2808_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x110y78     80'h00_0060_00_0000_0C08_FF2A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8167_4 ( .OUT(na8167_2), .IN1(na3290_1), .IN2(1'b1), .IN3(na4204_2), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x62y95     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8168_4 ( .OUT(na8168_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8168_5 ( .OUT(na8168_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8168_6 ( .RAM_O2(na8168_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8168_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y95     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8169_1 ( .OUT(na8169_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8169_2 ( .OUT(na8169_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8169_6 ( .RAM_O1(na8169_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8169_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y96     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8170_4 ( .OUT(na8170_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8170_5 ( .OUT(na8170_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8170_6 ( .RAM_O2(na8170_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8170_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y96     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8171_1 ( .OUT(na8171_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8171_2 ( .OUT(na8171_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8171_6 ( .RAM_O1(na8171_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8171_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y95     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8172_4 ( .OUT(na8172_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8172_5 ( .OUT(na8172_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8172_6 ( .RAM_O2(na8172_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8172_2_i), .COMP_OUT(1'b0) );
// C_AND////      x68y68     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8173_1 ( .OUT(na8173_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2554_1), .IN7(1'b1), .IN8(~na2556_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x76y72     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8174_4 ( .OUT(na8174_2), .IN1(na2566_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x70y74     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8175_1 ( .OUT(na8175_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2566_1), .IN6(1'b1), .IN7(na2558_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x58y85     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8176_1 ( .OUT(na8176_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2564_1), .IN7(1'b1), .IN8(na2556_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y59     80'h00_0018_00_0000_0C88_1CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8177_1 ( .OUT(na8177_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2557_1), .IN7(~na2558_1), .IN8(~na2556_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y95     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8178_1 ( .OUT(na8178_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8178_2 ( .OUT(na8178_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8178_6 ( .RAM_O1(na8178_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8178_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y94     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8179_4 ( .OUT(na8179_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8179_5 ( .OUT(na8179_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8179_6 ( .RAM_O2(na8179_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8179_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y94     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8180_1 ( .OUT(na8180_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8180_2 ( .OUT(na8180_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8180_6 ( .RAM_O1(na8180_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8180_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y93     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8181_4 ( .OUT(na8181_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8181_5 ( .OUT(na8181_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8181_6 ( .RAM_O2(na8181_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8181_2_i), .COMP_OUT(1'b0) );
// C_AND////      x89y102     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8182_1 ( .OUT(na8182_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na279_1), .IN6(na5452_1), .IN7(1'b1), .IN8(na272_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y76     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8183_1 ( .OUT(na8183_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3327_2), .IN6(na5953_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x51y78     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8184_4 ( .OUT(na8184_2), .IN1(~na3327_2), .IN2(na5953_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x114y69     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8185_4 ( .OUT(na8185_2), .IN1(na5218_1), .IN2(na9783_2), .IN3(na2163_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y66     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8186_1 ( .OUT(na8186_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3180_1), .IN6(1'b1), .IN7(na2163_1), .IN8(na5222_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y102     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8187_1 ( .OUT(na8187_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na279_1), .IN6(1'b1), .IN7(na5448_2), .IN8(na272_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y93     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8188_1 ( .OUT(na8188_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8188_2 ( .OUT(na8188_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8188_6 ( .RAM_O1(na8188_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8188_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y92     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8189_4 ( .OUT(na8189_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8189_5 ( .OUT(na8189_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8189_6 ( .RAM_O2(na8189_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8189_2_i), .COMP_OUT(1'b0) );
// C_///AND/      x95y110     80'h00_0060_00_0000_0C08_FF23
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8190_4 ( .OUT(na8190_2), .IN1(1'b1), .IN2(~na5223_2), .IN3(na3292_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y92     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8191_1 ( .OUT(na8191_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8191_2 ( .OUT(na8191_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8191_6 ( .RAM_O1(na8191_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8191_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x93y111     80'h00_0078_00_0000_0C88_2A2C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8192_1 ( .OUT(na8192_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3297_1), .IN6(1'b1), .IN7(na3357_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8192_4 ( .OUT(na8192_2), .IN1(1'b1), .IN2(na5223_2), .IN3(na3292_1), .IN4(~na6626_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y91     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8193_4 ( .OUT(na8193_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8193_5 ( .OUT(na8193_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8193_6 ( .RAM_O2(na8193_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8193_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y91     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8194_1 ( .OUT(na8194_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8194_2 ( .OUT(na8194_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8194_6 ( .RAM_O1(na8194_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8194_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y90     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8195_4 ( .OUT(na8195_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8195_5 ( .OUT(na8195_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8195_6 ( .RAM_O2(na8195_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8195_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y90     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8196_1 ( .OUT(na8196_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8196_2 ( .OUT(na8196_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8196_6 ( .RAM_O1(na8196_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8196_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x90y92     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8197_1 ( .OUT(na8197_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3354_1), .IN6(1'b1), .IN7(na3301_1), .IN8(~na6626_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y89     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8198_4 ( .OUT(na8198_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8198_5 ( .OUT(na8198_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8198_6 ( .RAM_O2(na8198_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8198_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y89     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8199_1 ( .OUT(na8199_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8199_2 ( .OUT(na8199_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8199_6 ( .RAM_O1(na8199_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8199_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y88     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8200_4 ( .OUT(na8200_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8200_5 ( .OUT(na8200_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8200_6 ( .RAM_O2(na8200_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8200_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y88     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8201_1 ( .OUT(na8201_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8201_2 ( .OUT(na8201_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8201_6 ( .RAM_O1(na8201_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8201_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y87     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8202_4 ( .OUT(na8202_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8202_5 ( .OUT(na8202_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8202_6 ( .RAM_O2(na8202_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8202_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y87     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8203_1 ( .OUT(na8203_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8203_2 ( .OUT(na8203_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8203_6 ( .RAM_O1(na8203_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8203_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y88     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8204_4 ( .OUT(na8204_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8204_5 ( .OUT(na8204_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8204_6 ( .RAM_O2(na8204_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8204_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y88     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8205_1 ( .OUT(na8205_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8205_2 ( .OUT(na8205_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8205_6 ( .RAM_O1(na8205_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8205_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y87     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8206_4 ( .OUT(na8206_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8206_5 ( .OUT(na8206_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8206_6 ( .RAM_O2(na8206_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8206_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y87     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8207_1 ( .OUT(na8207_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8207_2 ( .OUT(na8207_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8207_6 ( .RAM_O1(na8207_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8207_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y86     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8208_4 ( .OUT(na8208_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8208_5 ( .OUT(na8208_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8208_6 ( .RAM_O2(na8208_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8208_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y86     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8209_1 ( .OUT(na8209_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8209_2 ( .OUT(na8209_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8209_6 ( .RAM_O1(na8209_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8209_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y85     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8210_4 ( .OUT(na8210_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8210_5 ( .OUT(na8210_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8210_6 ( .RAM_O2(na8210_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8210_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y85     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8211_1 ( .OUT(na8211_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8211_2 ( .OUT(na8211_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8211_6 ( .RAM_O1(na8211_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8211_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y84     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8212_4 ( .OUT(na8212_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8212_5 ( .OUT(na8212_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8212_6 ( .RAM_O2(na8212_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8212_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y84     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8213_1 ( .OUT(na8213_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8213_2 ( .OUT(na8213_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8213_6 ( .RAM_O1(na8213_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8213_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y83     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8214_4 ( .OUT(na8214_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8214_5 ( .OUT(na8214_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8214_6 ( .RAM_O2(na8214_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8214_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y83     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8215_1 ( .OUT(na8215_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8215_2 ( .OUT(na8215_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8215_6 ( .RAM_O1(na8215_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8215_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y82     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8216_4 ( .OUT(na8216_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8216_5 ( .OUT(na8216_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8216_6 ( .RAM_O2(na8216_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8216_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y82     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8217_1 ( .OUT(na8217_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8217_2 ( .OUT(na8217_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8217_6 ( .RAM_O1(na8217_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8217_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y81     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8218_4 ( .OUT(na8218_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8218_5 ( .OUT(na8218_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8218_6 ( .RAM_O2(na8218_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8218_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y81     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8219_1 ( .OUT(na8219_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8219_2 ( .OUT(na8219_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6648_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8219_6 ( .RAM_O1(na8219_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8219_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y96     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8220_4 ( .OUT(na8220_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2882_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8220_6 ( .RAM_O2(na8220_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8220_2), .COMP_OUT(1'b0) );
// C_AND////      x61y96     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8221_1 ( .OUT(na8221_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2882_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8221_6 ( .RAM_O1(na8221_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8221_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y95     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8222_4 ( .OUT(na8222_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2882_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8222_6 ( .RAM_O2(na8222_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8222_2), .COMP_OUT(1'b0) );
// C_AND////      x61y95     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8223_1 ( .OUT(na8223_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2882_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8223_6 ( .RAM_O1(na8223_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8223_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y96     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8224_4 ( .OUT(na8224_2), .IN1(1'b1), .IN2(na2881_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8224_6 ( .RAM_O2(na8224_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8224_2), .COMP_OUT(1'b0) );
// C_AND////      x63y96     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8225_1 ( .OUT(na8225_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2881_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8225_6 ( .RAM_O1(na8225_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8225_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y95     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8226_4 ( .OUT(na8226_2), .IN1(1'b1), .IN2(na2881_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8226_6 ( .RAM_O2(na8226_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8226_2), .COMP_OUT(1'b0) );
// C_AND////      x63y95     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8227_1 ( .OUT(na8227_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2881_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8227_6 ( .RAM_O1(na8227_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8227_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y94     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8228_4 ( .OUT(na8228_2), .IN1(1'b1), .IN2(na2881_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8228_6 ( .RAM_O2(na8228_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8228_2), .COMP_OUT(1'b0) );
// C_AND////      x63y94     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8229_1 ( .OUT(na8229_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2881_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8229_6 ( .RAM_O1(na8229_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8229_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y93     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8230_4 ( .OUT(na8230_2), .IN1(1'b1), .IN2(na2881_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8230_6 ( .RAM_O2(na8230_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8230_2), .COMP_OUT(1'b0) );
// C_AND////      x63y93     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8231_1 ( .OUT(na8231_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2881_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8231_6 ( .RAM_O1(na8231_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8231_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y92     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8232_4 ( .OUT(na8232_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2880_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8232_6 ( .RAM_O2(na8232_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8232_2), .COMP_OUT(1'b0) );
// C_AND////      x63y92     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8233_1 ( .OUT(na8233_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2880_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8233_6 ( .RAM_O1(na8233_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8233_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y91     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8234_4 ( .OUT(na8234_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2880_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8234_6 ( .RAM_O2(na8234_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8234_2), .COMP_OUT(1'b0) );
// C_AND////      x63y91     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8235_1 ( .OUT(na8235_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2880_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8235_6 ( .RAM_O1(na8235_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8235_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y90     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8236_4 ( .OUT(na8236_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2880_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8236_6 ( .RAM_O2(na8236_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8236_2), .COMP_OUT(1'b0) );
// C_AND////      x63y90     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8237_1 ( .OUT(na8237_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2880_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8237_6 ( .RAM_O1(na8237_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8237_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y89     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8238_4 ( .OUT(na8238_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2880_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8238_6 ( .RAM_O2(na8238_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8238_2), .COMP_OUT(1'b0) );
// C_AND////      x63y89     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8239_1 ( .OUT(na8239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2880_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8239_6 ( .RAM_O1(na8239_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8239_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y88     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8240_4 ( .OUT(na8240_2), .IN1(na2888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8240_6 ( .RAM_O2(na8240_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8240_2), .COMP_OUT(1'b0) );
// C_AND////      x61y88     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8241_1 ( .OUT(na8241_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2888_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8241_6 ( .RAM_O1(na8241_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8241_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y87     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8242_4 ( .OUT(na8242_2), .IN1(na2888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8242_6 ( .RAM_O2(na8242_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8242_2), .COMP_OUT(1'b0) );
// C_AND////      x61y87     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8243_1 ( .OUT(na8243_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2888_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8243_6 ( .RAM_O1(na8243_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8243_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y88     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8244_4 ( .OUT(na8244_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2887_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8244_6 ( .RAM_O2(na8244_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8244_2), .COMP_OUT(1'b0) );
// C_AND////      x63y88     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8245_1 ( .OUT(na8245_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2887_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8245_6 ( .RAM_O1(na8245_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8245_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y87     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8246_4 ( .OUT(na8246_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2887_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8246_6 ( .RAM_O2(na8246_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8246_2), .COMP_OUT(1'b0) );
// C_AND////      x63y87     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8247_1 ( .OUT(na8247_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2887_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8247_6 ( .RAM_O1(na8247_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8247_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y86     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8248_4 ( .OUT(na8248_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2887_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8248_6 ( .RAM_O2(na8248_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8248_2), .COMP_OUT(1'b0) );
// C_AND////      x63y86     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8249_1 ( .OUT(na8249_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2887_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8249_6 ( .RAM_O1(na8249_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8249_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y85     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8250_4 ( .OUT(na8250_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2887_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8250_6 ( .RAM_O2(na8250_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8250_2), .COMP_OUT(1'b0) );
// C_AND////      x63y85     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8251_1 ( .OUT(na8251_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2887_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8251_6 ( .RAM_O1(na8251_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8251_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y84     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8252_4 ( .OUT(na8252_2), .IN1(1'b1), .IN2(na2886_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8252_6 ( .RAM_O2(na8252_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8252_2), .COMP_OUT(1'b0) );
// C_AND////      x63y84     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8253_1 ( .OUT(na8253_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2886_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8253_6 ( .RAM_O1(na8253_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8253_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y83     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8254_4 ( .OUT(na8254_2), .IN1(1'b1), .IN2(na2886_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8254_6 ( .RAM_O2(na8254_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8254_2), .COMP_OUT(1'b0) );
// C_AND////      x63y83     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8255_1 ( .OUT(na8255_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2886_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8255_6 ( .RAM_O1(na8255_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8255_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y82     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8256_4 ( .OUT(na8256_2), .IN1(1'b1), .IN2(na2886_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8256_6 ( .RAM_O2(na8256_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8256_2), .COMP_OUT(1'b0) );
// C_AND////      x63y82     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8257_1 ( .OUT(na8257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2886_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8257_6 ( .RAM_O1(na8257_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8257_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y81     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8258_4 ( .OUT(na8258_2), .IN1(1'b1), .IN2(na2886_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8258_6 ( .RAM_O2(na8258_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8258_2), .COMP_OUT(1'b0) );
// C_AND////      x63y81     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8259_1 ( .OUT(na8259_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2886_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8259_6 ( .RAM_O1(na8259_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8259_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x35y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8260_1 ( .OUT(na8260_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8260_6 ( .RAM_O1(na8260_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8260_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x35y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8261_1 ( .OUT(na8261_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8261_6 ( .RAM_O1(na8261_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8261_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y57     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8262_4 ( .OUT(na8262_2), .IN1(1'b1), .IN2(na3229_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8262_6 ( .RAM_O2(na8262_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8262_2), .COMP_OUT(1'b0) );
// C_///AND/      x27y49     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8263_4 ( .OUT(na8263_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2892_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8263_6 ( .RAM_O2(na8263_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8263_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y56     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8264_4 ( .OUT(na8264_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8264_6 ( .RAM_O2(na8264_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8264_2), .COMP_OUT(1'b0) );
// C_AND////      x28y56     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8265_1 ( .OUT(na8265_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8265_6 ( .RAM_O1(na8265_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8265_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y55     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8266_4 ( .OUT(na8266_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8266_6 ( .RAM_O2(na8266_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8266_2), .COMP_OUT(1'b0) );
// C_ORAND////      x83y78     80'h00_0018_00_0000_0888_DD77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8267_1 ( .OUT(na8267_1), .IN1(~na88_1), .IN2(~na9171_2), .IN3(~na63_1), .IN4(~na9175_2), .IN5(~na95_1), .IN6(na15_1), .IN7(~na97_2),
                      .IN8(na9141_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y55     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8268_1 ( .OUT(na8268_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8268_6 ( .RAM_O1(na8268_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8268_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y54     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8269_4 ( .OUT(na8269_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8269_6 ( .RAM_O2(na8269_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8269_2), .COMP_OUT(1'b0) );
// C_AND////      x28y54     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8270_1 ( .OUT(na8270_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8270_6 ( .RAM_O1(na8270_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8270_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x95y94     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8271_1 ( .OUT(na8271_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na104_1), .IN7(~na2937_2), .IN8(na6692_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y89     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a8272_1 ( .OUT(na8272_1), .IN1(1'b1), .IN2(1'b1), .IN3(na2937_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na2971_1), .IN7(1'b0), .IN8(~na2976_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y53     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8273_4 ( .OUT(na8273_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8273_6 ( .RAM_O2(na8273_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8273_2), .COMP_OUT(1'b0) );
// C_///ORAND/      x95y100     80'h00_0060_00_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a8274_4 ( .OUT(na8274_2), .IN1(na8272_1), .IN2(~na2935_1), .IN3(na128_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y47     80'h00_0078_00_0000_0C66_3C90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8275_1 ( .OUT(na8275_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na5687_1), .IN7(1'b0), .IN8(~na2590_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8275_4 ( .OUT(na8275_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5688_1), .IN4(~na2592_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y53     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8276_1 ( .OUT(na8276_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8276_6 ( .RAM_O1(na8276_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8276_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x58y50     80'h00_0078_00_0000_0C66_AA5A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8277_1 ( .OUT(na8277_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2584_2), .IN6(1'b0), .IN7(na5684_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8277_4 ( .OUT(na8277_2), .IN1(na5686_1), .IN2(1'b0), .IN3(~na2588_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x56y38     80'h00_0078_00_0000_0C66_3C90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8278_1 ( .OUT(na8278_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na5687_1), .IN7(1'b0), .IN8(~na2580_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8278_4 ( .OUT(na8278_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5688_1), .IN4(~na2582_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y52     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8279_4 ( .OUT(na8279_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8279_6 ( .RAM_O2(na8279_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8279_2), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x55y38     80'h00_0078_00_0000_0C66_AA09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8280_1 ( .OUT(na8280_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2574_2), .IN6(1'b0), .IN7(na5684_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8280_4 ( .OUT(na8280_2), .IN1(na5686_1), .IN2(~na2578_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8281_1 ( .OUT(na8281_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8281_6 ( .RAM_O1(na8281_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8281_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y51     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8282_4 ( .OUT(na8282_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8282_6 ( .RAM_O2(na8282_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8282_2), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x66y54     80'h00_0078_00_0000_0C66_3A09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8283_1 ( .OUT(na8283_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2576_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na5962_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8283_4 ( .OUT(na8283_2), .IN1(na2574_2), .IN2(~na5948_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y51     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8284_1 ( .OUT(na8284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8284_6 ( .RAM_O1(na8284_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8284_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x62y51     80'h00_0078_00_0000_0C66_9009
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8285_1 ( .OUT(na8285_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na5964_2), .IN8(na2580_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8285_4 ( .OUT(na8285_2), .IN1(~na5963_2), .IN2(na2578_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x79y59     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8286_4 ( .OUT(na8286_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na5965_2), .IN4(na2582_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x56y37     80'h00_0078_00_0000_0C66_5AC3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8287_1 ( .OUT(na8287_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2574_2), .IN6(1'b0), .IN7(~na5684_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8287_4 ( .OUT(na8287_2), .IN1(1'b0), .IN2(~na5687_2), .IN3(1'b0), .IN4(na2580_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x56y42     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8288_1 ( .OUT(na8288_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2576_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na5685_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y40     80'h00_0078_00_0000_0C66_0990
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8289_1 ( .OUT(na8289_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na5686_2), .IN6(na2578_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8289_4 ( .OUT(na8289_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na5688_2), .IN4(na2582_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8290_4 ( .OUT(na8290_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8290_6 ( .RAM_O2(na8290_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8290_2), .COMP_OUT(1'b0) );
// C_AND////      x28y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8291_1 ( .OUT(na8291_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8291_6 ( .RAM_O1(na8291_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8291_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x61y44     80'h00_0078_00_0000_0C66_90A5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8292_1 ( .OUT(na8292_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5932_2), .IN8(~na2580_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8292_4 ( .OUT(na8292_2), .IN1(~na2576_2), .IN2(1'b0), .IN3(na5932_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8293_4 ( .OUT(na8293_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8293_6 ( .RAM_O2(na8293_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8293_2), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x58y46     80'h00_0078_00_0000_0C66_093A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8294_1 ( .OUT(na8294_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5935_2), .IN6(~na2578_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8294_4 ( .OUT(na8294_2), .IN1(na5935_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na2582_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x57y48     80'h00_0078_00_0000_0C66_5A90
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8295_1 ( .OUT(na8295_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2584_2), .IN6(1'b0), .IN7(~na5684_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8295_4 ( .OUT(na8295_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na5688_2), .IN4(na2592_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x75y61     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8296_4 ( .OUT(na8296_2), .IN1(1'b0), .IN2(na2586_2), .IN3(1'b0), .IN4(~na5685_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x58y48     80'h00_0078_00_0000_0C66_A5C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8297_1 ( .OUT(na8297_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na5686_2), .IN6(1'b0), .IN7(na2588_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8297_4 ( .OUT(na8297_2), .IN1(1'b0), .IN2(~na5687_2), .IN3(1'b0), .IN4(na2590_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8298_1 ( .OUT(na8298_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8298_6 ( .RAM_O1(na8298_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8298_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y64     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8299_4 ( .OUT(na8299_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8299_6 ( .RAM_O2(na8299_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8299_2), .COMP_OUT(1'b0) );
// C_OR////      x58y52     80'h00_0018_00_0000_0EEE_3777
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8300_1 ( .OUT(na8300_1), .IN1(~na1372_1), .IN2(~na8295_2), .IN3(~na1387_2), .IN4(~na8297_2), .IN5(~na8296_2), .IN6(~na8295_1),
                      .IN7(1'b0), .IN8(~na8297_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y64     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8301_1 ( .OUT(na8301_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8301_6 ( .RAM_O1(na8301_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8301_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x66y64     80'h00_0078_00_0000_0C66_C55A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8302_1 ( .OUT(na8302_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na2584_2), .IN6(1'b0), .IN7(1'b0), .IN8(na5931_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8302_4 ( .OUT(na8302_2), .IN1(na5935_2), .IN2(1'b0), .IN3(~na2588_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y63     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8303_4 ( .OUT(na8303_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8303_6 ( .RAM_O2(na8303_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8303_2), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x66y63     80'h00_0078_00_0000_0C66_90A3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8304_1 ( .OUT(na8304_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5932_2), .IN8(~na2590_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8304_4 ( .OUT(na8304_2), .IN1(1'b0), .IN2(~na2586_2), .IN3(na5932_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x63y53     80'h00_0018_00_0000_0C66_3A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8305_1 ( .OUT(na8305_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5935_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na2592_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y63     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8306_1 ( .OUT(na8306_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8306_6 ( .RAM_O1(na8306_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8306_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x77y73     80'h00_0078_00_0000_0C66_3C09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8307_1 ( .OUT(na8307_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2586_2), .IN7(1'b0), .IN8(~na5962_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8307_4 ( .OUT(na8307_2), .IN1(na2584_2), .IN2(~na5948_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y62     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8308_4 ( .OUT(na8308_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8308_6 ( .RAM_O2(na8308_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8308_2), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x74y70     80'h00_0078_00_0000_0C66_90A5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8309_1 ( .OUT(na8309_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na5964_2), .IN8(na2590_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8309_4 ( .OUT(na8309_2), .IN1(~na5963_2), .IN2(1'b0), .IN3(na2588_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x75y62     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8310_4 ( .OUT(na8310_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na5965_2), .IN4(na2592_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y62     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8311_1 ( .OUT(na8311_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8311_6 ( .RAM_O1(na8311_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8311_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x80y75     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8312_1 ( .OUT(na8312_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na380_2), .IN8(na2572_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y60     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8313_4 ( .OUT(na8313_2), .IN1(na2566_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na9623_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y75     80'h00_0018_00_0000_0888_5111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8314_1 ( .OUT(na8314_1), .IN1(~na2570_1), .IN2(~na2571_1), .IN3(~na2568_1), .IN4(~na2573_1), .IN5(~na2569_1), .IN6(~na2567_1),
                      .IN7(~na2558_1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y76     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8315_4 ( .OUT(na8315_2), .IN1(1'b1), .IN2(na2557_1), .IN3(1'b1), .IN4(~na2556_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y61     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8316_4 ( .OUT(na8316_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8316_6 ( .RAM_O2(na8316_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8316_2), .COMP_OUT(1'b0) );
// C_ORAND////      x77y69     80'h00_0018_00_0000_0888_ECC5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8317_1 ( .OUT(na8317_1), .IN1(~na2555_1), .IN2(1'b0), .IN3(1'b0), .IN4(na3532_1), .IN5(1'b0), .IN6(na9210_2), .IN7(na380_2),
                      .IN8(na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x76y68     80'h00_0018_00_0000_0C88_31FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8318_1 ( .OUT(na8318_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2566_1), .IN6(~na2557_1), .IN7(1'b1), .IN8(~na9623_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x78y74     80'h00_0018_00_0000_0EEE_C537
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8319_1 ( .OUT(na8319_1), .IN1(~na3535_1), .IN2(~na2554_1), .IN3(1'b0), .IN4(~na393_2), .IN5(~na2555_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na2556_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y61     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8320_1 ( .OUT(na8320_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8320_6 ( .RAM_O1(na8320_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8320_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y60     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8321_4 ( .OUT(na8321_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8321_6 ( .RAM_O2(na8321_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8321_2), .COMP_OUT(1'b0) );
// C_///AND/      x82y84     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8322_4 ( .OUT(na8322_2), .IN1(na3305_1), .IN2(1'b1), .IN3(na561_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x68y118     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8323_1 ( .OUT(na8323_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1388_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na3309_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y112     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8324_4 ( .OUT(na8324_2), .IN1(1'b1), .IN2(na3317_1), .IN3(1'b1), .IN4(na1407_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x126y68     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a8325_4 ( .OUT(na8325_2), .IN1(1'b0), .IN2(na647_1), .IN3(na9180_2), .IN4(na154_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8326_1 ( .OUT(na8326_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8326_6 ( .RAM_O1(na8326_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8326_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x109y78     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8327_1 ( .OUT(na8327_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na212_1), .IN6(na2935_1), .IN7(na2937_2), .IN8(na174_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x110y67     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8328_4 ( .OUT(na8328_2), .IN1(1'b1), .IN2(na99_2), .IN3(1'b1), .IN4(~na194_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x132y78     80'h00_0018_00_0040_0C94_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a8329_1 ( .OUT(na8329_1), .IN1(1'b1), .IN2(1'b0), .IN3(na3544_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2894_2), .IN7(1'b1), .IN8(~na3543_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x112y73     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8330_1 ( .OUT(na8330_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na6485_1), .IN6(~na9830_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y59     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8331_4 ( .OUT(na8331_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8331_6 ( .RAM_O2(na8331_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8331_2), .COMP_OUT(1'b0) );
// C_///AND/      x93y91     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8332_4 ( .OUT(na8332_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na3276_1), .IN4(~na6497_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y94     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8333_1 ( .OUT(na8333_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3549_1), .IN7(~na3301_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8334_1 ( .OUT(na8334_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8334_6 ( .RAM_O1(na8334_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8334_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8335_4 ( .OUT(na8335_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8335_6 ( .RAM_O2(na8335_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8335_2), .COMP_OUT(1'b0) );
// C_AND////      x28y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8336_1 ( .OUT(na8336_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8336_6 ( .RAM_O1(na8336_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8336_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x123y69     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a8337_4 ( .OUT(na8337_2), .IN1(~na488_1), .IN2(~na981_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y67     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8338_1 ( .OUT(na8338_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na430_1), .IN8(~na3552_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x110y65     80'h00_0018_00_0000_0EEE_E5D3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8339_1 ( .OUT(na8339_1), .IN1(1'b0), .IN2(~na9955_2), .IN3(~na7311_1), .IN4(na7310_1), .IN5(~na8337_2), .IN6(1'b0), .IN7(na8338_1),
                      .IN8(na7312_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8340_4 ( .OUT(na8340_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8340_6 ( .RAM_O2(na8340_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8340_2), .COMP_OUT(1'b0) );
// C_AND////      x118y69     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8341_1 ( .OUT(na8341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na3219_2), .IN8(na3227_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8342_1 ( .OUT(na8342_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8342_6 ( .RAM_O1(na8342_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8342_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x37y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8343_1 ( .OUT(na8343_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8343_6 ( .RAM_O1(na8343_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8343_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x86y78     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8344_1 ( .OUT(na8344_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1524_1), .IN7(na1248_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y64     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a8345_1 ( .OUT(na8345_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1132_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1595_2), .IN7(1'b0), .IN8(~na1531_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x90y72     80'h00_0018_00_0000_0EEE_7BDA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8346_1 ( .OUT(na8346_1), .IN1(na7362_2), .IN2(1'b0), .IN3(~na7359_1), .IN4(na8344_1), .IN5(na7360_1), .IN6(~na8345_1), .IN7(~na7359_2),
                      .IN8(~na7361_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y51     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8347_1 ( .OUT(na8347_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8347_6 ( .RAM_O1(na8347_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8347_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x52y72     80'h00_0018_00_0000_0888_8828
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8348_1 ( .OUT(na8348_1), .IN1(na2342_1), .IN2(na2367_1), .IN3(na2306_1), .IN4(~na5955_2), .IN5(na2334_1), .IN6(na2325_1),
                      .IN7(na2380_1), .IN8(na2337_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x76y90     80'h00_0060_00_0000_0C06_FF36
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8349_4 ( .OUT(na8349_2), .IN1(na2389_1), .IN2(na5953_1), .IN3(1'b0), .IN4(~na8348_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8350_4 ( .OUT(na8350_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8350_6 ( .RAM_O2(na8350_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8350_2), .COMP_OUT(1'b0) );
// C_AND////      x37y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8351_1 ( .OUT(na8351_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8351_6 ( .RAM_O1(na8351_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8351_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x89y92     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8352_1 ( .OUT(na8352_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3588_1), .IN6(~na3213_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8353_4 ( .OUT(na8353_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8353_6 ( .RAM_O2(na8353_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8353_2), .COMP_OUT(1'b0) );
// C_AND////      x37y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8354_1 ( .OUT(na8354_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8354_6 ( .RAM_O1(na8354_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8354_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///XOR/      x130y115     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8355_4 ( .OUT(na8355_2), .IN1(na6055_1), .IN2(~na318_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8356_1 ( .OUT(na8356_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8356_6 ( .RAM_O1(na8356_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8356_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x129y115     80'h00_0078_00_0000_0C66_CA5A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8357_1 ( .OUT(na8357_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na6055_2), .IN6(1'b0), .IN7(1'b0), .IN8(na321_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8357_4 ( .OUT(na8357_2), .IN1(na6055_1), .IN2(1'b0), .IN3(~na320_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x119y107     80'h00_0060_00_0000_0C08_FFC8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8358_4 ( .OUT(na8358_2), .IN1(na2733_1), .IN2(na3592_1), .IN3(1'b1), .IN4(na3665_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8359_1 ( .OUT(na8359_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8359_6 ( .RAM_O1(na8359_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8359_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x119y72     80'h00_0018_00_0000_0888_88CF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8360_1 ( .OUT(na8360_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1333_1), .IN5(na900_1), .IN6(na3345_1), .IN7(na1119_1),
                      .IN8(na3590_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y58     80'h00_0060_00_0000_0C08_FFC4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8361_4 ( .OUT(na8361_2), .IN1(~na2566_1), .IN2(na2557_1), .IN3(1'b1), .IN4(na2572_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x79y73     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a8362_4 ( .OUT(na8362_2), .IN1(~na3597_1), .IN2(~na9615_2), .IN3(~na2558_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x76y72     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8363_1 ( .OUT(na8363_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2565_1), .IN6(na8361_2), .IN7(1'b0), .IN8(na2556_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8364_4 ( .OUT(na8364_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8364_6 ( .RAM_O2(na8364_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8364_2), .COMP_OUT(1'b0) );
// C_///OR/      x73y62     80'h00_0060_00_0000_0C0E_FFBD
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a8365_4 ( .OUT(na8365_2), .IN1(~na3501_1), .IN2(na3525_1), .IN3(na3521_1), .IN4(~na8300_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8366_1 ( .OUT(na8366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8366_6 ( .RAM_O1(na8366_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8366_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x75y73     80'h00_0018_00_0000_0888_F37C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8367_1 ( .OUT(na8367_1), .IN1(1'b0), .IN2(na8365_2), .IN3(~na2558_1), .IN4(~na2556_1), .IN5(1'b0), .IN6(~na369_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8368_4 ( .OUT(na8368_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8368_6 ( .RAM_O2(na8368_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8368_2), .COMP_OUT(1'b0) );
// C_AND////      x37y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8369_1 ( .OUT(na8369_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8369_6 ( .RAM_O1(na8369_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8369_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x71y64     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8370_1 ( .OUT(na8370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2555_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na2556_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x74y97     80'h00_0078_00_0000_0CEE_5CD5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a8371_1 ( .OUT(na8371_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na8372_2), .IN7(~na1492_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a8371_4 ( .OUT(na8371_2), .IN1(~na1372_1), .IN2(1'b0), .IN3(~na9904_2), .IN4(na5435_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x75y92     80'h00_0060_00_0000_0C08_FF51
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8372_4 ( .OUT(na8372_2), .IN1(~na8367_1), .IN2(~na521_1), .IN3(~na3603_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x80y96     80'h00_0078_00_0000_0C88_3AC4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8373_1 ( .OUT(na8373_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2570_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na389_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8373_4 ( .OUT(na8373_2), .IN1(~na2584_2), .IN2(na2586_2), .IN3(1'b1), .IN4(na389_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x30y64     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8374_4 ( .OUT(na8374_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8374_5 ( .OUT(na8374_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8374_6 ( .RAM_O2(na8374_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8374_2_i), .COMP_OUT(1'b0) );
// C_AND///AND/      x81y86     80'h00_0078_00_0000_0C88_F15A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8375_1 ( .OUT(na8375_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2570_1), .IN6(~na387_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8375_4 ( .OUT(na8375_2), .IN1(na2570_1), .IN2(1'b1), .IN3(~na3307_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x30y64     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8376_1 ( .OUT(na8376_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8376_2 ( .OUT(na8376_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8376_6 ( .RAM_O1(na8376_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8376_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x87y64     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8377_4 ( .OUT(na8377_2), .IN1(~na2566_1), .IN2(~na2564_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y63     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8378_1 ( .OUT(na8378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2557_1), .IN7(1'b1), .IN8(~na3608_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y72     80'h00_0018_00_0000_0888_C573
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8379_1 ( .OUT(na8379_1), .IN1(1'b0), .IN2(~na2554_1), .IN3(~na3612_1), .IN4(~na3526_1), .IN5(~na2555_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na393_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x30y63     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8380_4 ( .OUT(na8380_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8380_5 ( .OUT(na8380_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8380_6 ( .RAM_O2(na8380_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8380_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x30y63     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8381_1 ( .OUT(na8381_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8381_2 ( .OUT(na8381_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8381_6 ( .RAM_O1(na8381_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8381_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x80y71     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8382_1 ( .OUT(na8382_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na3529_1), .IN7(1'b1), .IN8(~na3611_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND*/      x128y106     80'h00_0060_00_0000_0C07_FFF0
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a8383_4 ( .OUT(na8383_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND//O_0/AND/      x128y107     80'h00_0078_09_6000_FC88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8384_1 ( .OUT(na8384_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2796_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a8384_3 ( .COMP_OUT(na8384_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8384_4 ( .OUT(na8384_2), .IN1(1'b1), .IN2(na2795_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a8384_6 ( .COUTX(na8384_3), .POUTX(na8384_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8384_1), .OUT2(na8384_2), .COMP_OUT(na8384_3_i) );
// C_AND*//O_0/AND*/      x128y108     80'h00_0078_09_6000_F387_FAFA
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a8385_1 ( .OUT(na8385_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2793_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a8385_3 ( .COMP_OUT(na8385_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a8385_4 ( .OUT(na8385_2), .IN1(na2794_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a8385_6 ( .COUTX(na8385_3), .POUTX(na8385_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8385_1), .OUT2(na8385_2), .COMP_OUT(na8385_3_i) );
// C_AND//O_0/AND/      x128y109     80'h00_0078_09_6000_FC88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8386_1 ( .OUT(na8386_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2792_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a8386_3 ( .COMP_OUT(na8386_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8386_4 ( .OUT(na8386_2), .IN1(na2741_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a8386_6 ( .COUTX(na8386_3), .POUTX(na8386_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8386_1), .OUT2(na8386_2), .COMP_OUT(na8386_3_i) );
// C_AND*//O_0/AND*/      x128y110     80'h00_0078_09_6000_F387_CFFA
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a8387_1 ( .OUT(na8387_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2791_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a8387_3 ( .COMP_OUT(na8387_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a8387_4 ( .OUT(na8387_2), .IN1(na2790_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a8387_6 ( .COUTX(na8387_3), .POUTX(na8387_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8387_1), .OUT2(na8387_2), .COMP_OUT(na8387_3_i) );
// C_AND//O_0/AND/      x128y111     80'h00_0078_09_6000_FC88_F0F0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8388_1 ( .OUT(na8388_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a8388_3 ( .COMP_OUT(na8388_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8388_4 ( .OUT(na8388_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a8388_6 ( .COUTX(na8388_3), .POUTX(na8388_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8388_1), .OUT2(na8388_2), .COMP_OUT(na8388_3_i) );
// C_AND*//O_0/AND*/      x128y112     80'h00_0078_09_6000_F387_F0F0
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a8389_1 ( .OUT(na8389_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a8389_3 ( .COMP_OUT(na8389_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a8389_4 ( .OUT(na8389_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a8389_6 ( .COUTX(na8389_3), .POUTX(na8389_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8389_1), .OUT2(na8389_2), .COMP_OUT(na8389_3_i) );
// C_AND///AND/      x129y103     80'h00_0078_12_0000_0C88_F3FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8390_1 ( .OUT(na8390_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2933_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8390_4 ( .OUT(na8390_2), .IN1(1'b1), .IN2(na2933_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a8390_6 ( .COUTY1(na8390_4), .POUTY1(na8390_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8390_1), .OUT2(na8390_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x129y104     80'h00_0018_04_2056_5888_0CC0
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a8391_1 ( .OUT(na8391_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na8390_4), .PINX(1'b0), .PINY1(na8390_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a8391_3 ( .COMP_OUT(na8391_3_i), .COMB1(na8391_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a8391_6 ( .COUTY1(na8391_4), .COUTY2(na8391_5), .POUTY1(na8391_7), .CINX(1'b0), .CINY1(na8390_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na8390_7), .PINY2(1'b0), .OUT1(na8391_1), .OUT2(1'b0), .COMP_OUT(na8391_3_i) );
// C_MULTFa//O_O2//      x129y105     80'h00_0018_13_A477_34A6_0C0C
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a8392_1 ( .COUTX(na8392_3), .COUTY1(na8392_4), .COUTY2(na8392_5), .POUTY1(na8392_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na8391_4),
                      .CINY2(na8391_5), .PINX(1'b0), .PINY1(na8391_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x129y106     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a8393_1 ( .OUT(na8393_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na8392_4), .PINX(1'b0), .PINY1(na8392_7) );
C_O_0      #(.CPE_CFG ()) 
           _a8393_3 ( .COMP_OUT(na8393_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a8393_4 ( .OUT(na8393_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na8392_4), .PINX(1'b0), .PINY1(na8392_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a8393_6 ( .COUTX(na8393_3), .COUTY1(na8393_4), .COUTY2(na8393_5), .POUTY1(na8393_7), .POUTY2(na8393_8), .CINX(1'b0), .CINY1(na8392_4),
                      .CINY2(na8392_5), .PINX(1'b0), .PINY1(na8392_7), .PINY2(1'b0), .OUT1(na8393_1), .OUT2(na8393_2), .COMP_OUT(na8393_3_i) );
// C_MULT///MULT/      x129y107     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8394_1 ( .OUT1(na8394_1), .OUT2(na8394_2), .COUTY1(na8394_4), .COUTY2(na8394_5), .POUTY1(na8394_7), .POUTY2(na8394_8), .IN1(na8384_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8384_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8383_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(1'b0), .CINY1(na8393_4), .CINY2(na8393_5), .PINX(1'b0), .PINY1(na8393_7), .PINY2(na8393_8), .RAM_I1(1'b0),
                      .RAM_I2(1'b0) );
// C_MULT///MULT/      x129y108     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8395_1 ( .COUTX(na8395_3), .COUTY1(na8395_4), .COUTY2(na8395_5), .POUTX(na8395_6), .POUTY1(na8395_7), .POUTY2(na8395_8),
                      .IN1(~na8385_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na8385_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8384_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na8394_4), .CINY2(na8394_5), .PINX(1'b0), .PINY1(na8394_7), .PINY2(na8394_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x129y109     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8396_1 ( .COUTX(na8396_3), .COUTY1(na8396_4), .COUTY2(na8396_5), .POUTX(na8396_6), .POUTY1(na8396_7), .POUTY2(na8396_8),
                      .IN1(na8386_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8386_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8385_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na8395_4), .CINY2(na8395_5), .PINX(1'b0), .PINY1(na8395_7), .PINY2(na8395_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x129y110     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8397_1 ( .COUTX(na8397_3), .COUTY1(na8397_4), .COUTY2(na8397_5), .POUTX(na8397_6), .POUTY1(na8397_7), .POUTY2(na8397_8),
                      .IN1(~na8387_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na8387_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8386_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na8396_4), .CINY2(na8396_5), .PINX(1'b0), .PINY1(na8396_7), .PINY2(na8396_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x129y111     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8398_1 ( .COUTX(na8398_3), .COUTY1(na8398_4), .COUTY2(na8398_5), .POUTX(na8398_6), .POUTY1(na8398_7), .POUTY2(na8398_8),
                      .IN1(na8388_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8388_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8387_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na8397_4), .CINY2(na8397_5), .PINX(1'b0), .PINY1(na8397_7), .PINY2(na8397_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x129y112     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a8399_1 ( .COUTX(na8399_3), .COUTY1(na8399_4), .COUTY2(na8399_5), .POUTX(na8399_6), .POUTY1(na8399_7), .POUTY2(na8399_8),
                      .IN1(~na8389_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na8389_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8388_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na8398_4), .CINY2(na8398_5), .PINX(1'b0), .PINY1(na8398_7), .PINY2(na8398_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x129y113     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a8400_3 ( .COMP_OUT(na8400_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a8400_4 ( .OUT(na8400_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na8399_4), .PINX(1'b0), .PINY1(na8399_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a8400_6 ( .COUTX(na8400_3), .POUTX(na8400_6), .CINX(1'b0), .CINY1(na8399_4), .CINY2(na8399_5), .PINX(1'b0), .PINY1(na8399_7),
                      .PINY2(na8399_8), .OUT1(1'b0), .OUT2(na8400_2), .COMP_OUT(na8400_3_i) );
// C_AND///AND/      x130y104     80'h00_0078_12_0000_0C88_F0F0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8401_1 ( .OUT(na8401_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8401_4 ( .OUT(na8401_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a8401_6 ( .COUTY1(na8401_4), .POUTY1(na8401_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8401_1), .OUT2(na8401_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x130y105     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a8402_1 ( .OUT(na8402_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na8392_3), .CINY1(na8401_4), .PINX(1'b0), .PINY1(na8401_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a8402_3 ( .COMP_OUT(na8402_3_i), .COMB1(na8402_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a8402_6 ( .COUTY1(na8402_4), .COUTY2(na8402_5), .POUTY1(na8402_7), .CINX(na8392_3), .CINY1(na8401_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na8401_7), .PINY2(1'b0), .OUT1(na8402_1), .OUT2(1'b0), .COMP_OUT(na8402_3_i) );
// C_MULTFb//O_O2//      x130y106     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a8403_1 ( .COUTX(na8403_3), .COUTY1(na8403_4), .COUTY2(na8403_5), .POUTY1(na8403_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na8393_3), .CINY1(na8402_4),
                      .CINY2(na8402_5), .PINX(1'b0), .PINY1(na8402_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x130y107     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a8404_1 ( .OUT(na8404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na8403_4), .PINX(1'b0), .PINY1(na8403_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a8404_3 ( .COMP_OUT(na8404_3_i), .COMB1(1'b0), .COMB2(na8404_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a8404_4 ( .OUT(na8404_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na8403_4), .PINX(1'b0), .PINY1(na8403_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a8404_6 ( .COUTX(na8404_3), .COUTY1(na8404_4), .COUTY2(na8404_5), .POUTY1(na8404_7), .POUTY2(na8404_8), .CINX(1'b0), .CINY1(na8403_4),
                      .CINY2(na8403_5), .PINX(1'b0), .PINY1(na8403_7), .PINY2(1'b0), .OUT1(na8404_1), .OUT2(na8404_2), .COMP_OUT(na8404_3_i) );
// C_MULT///MULT/      x130y108     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8405_1 ( .OUT1(na8405_1), .OUT2(na8405_2), .COUTY1(na8405_4), .COUTY2(na8405_5), .POUTY1(na8405_7), .POUTY2(na8405_8), .IN1(~na8384_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na8384_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8383_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na8395_3), .CINY1(na8404_4), .CINY2(na8404_5), .PINX(na8395_6), .PINY1(na8404_7), .PINY2(na8404_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x130y109     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8406_1 ( .COUTX(na8406_3), .COUTY1(na8406_4), .COUTY2(na8406_5), .POUTX(na8406_6), .POUTY1(na8406_7), .POUTY2(na8406_8),
                      .IN1(na8385_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8385_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8384_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na8396_3), .CINY1(na8405_4), .CINY2(na8405_5), .PINX(na8396_6), .PINY1(na8405_7), .PINY2(na8405_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x130y110     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8407_1 ( .COUTX(na8407_3), .COUTY1(na8407_4), .COUTY2(na8407_5), .POUTX(na8407_6), .POUTY1(na8407_7), .POUTY2(na8407_8),
                      .IN1(~na8386_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na8386_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8385_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na8397_3), .CINY1(na8406_4), .CINY2(na8406_5), .PINX(na8397_6), .PINY1(na8406_7), .PINY2(na8406_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x130y111     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8408_1 ( .COUTX(na8408_3), .COUTY1(na8408_4), .COUTY2(na8408_5), .POUTX(na8408_6), .POUTY1(na8408_7), .POUTY2(na8408_8),
                      .IN1(na8387_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8387_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8386_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na8398_3), .CINY1(na8407_4), .CINY2(na8407_5), .PINX(na8398_6), .PINY1(na8407_7), .PINY2(na8407_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x130y112     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8409_1 ( .COUTX(na8409_3), .COUTY1(na8409_4), .COUTY2(na8409_5), .POUTX(na8409_6), .POUTY1(na8409_7), .POUTY2(na8409_8),
                      .IN1(~na8388_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na8388_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8387_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na8399_3), .CINY1(na8408_4), .CINY2(na8408_5), .PINX(na8399_6), .PINY1(na8408_7), .PINY2(na8408_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x130y113     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a8410_1 ( .COUTX(na8410_3), .COUTY1(na8410_4), .COUTY2(na8410_5), .POUTX(na8410_6), .POUTY1(na8410_7), .POUTY2(na8410_8),
                      .IN1(na8389_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8389_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8388_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na8400_3), .CINY1(na8409_4), .CINY2(na8409_5), .PINX(na8400_6), .PINY1(na8409_7), .PINY2(na8409_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x130y114     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a8411_3 ( .COMP_OUT(na8411_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a8411_4 ( .OUT(na8411_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na8410_4), .PINX(1'b0), .PINY1(na8410_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a8411_6 ( .COUTX(na8411_3), .POUTX(na8411_6), .CINX(1'b0), .CINY1(na8410_4), .CINY2(na8410_5), .PINX(1'b0), .PINY1(na8410_7),
                      .PINY2(na8410_8), .OUT1(1'b0), .OUT2(na8411_2), .COMP_OUT(na8411_3_i) );
// C_AND///AND/      x131y105     80'h00_0078_12_0000_0C88_F0F0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8412_1 ( .OUT(na8412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8412_4 ( .OUT(na8412_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a8412_6 ( .COUTY1(na8412_4), .POUTY1(na8412_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na8412_1), .OUT2(na8412_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x131y106     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a8413_1 ( .OUT(na8413_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na8403_3), .CINY1(na8412_4), .PINX(1'b0), .PINY1(na8412_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a8413_3 ( .COMP_OUT(na8413_3_i), .COMB1(na8413_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a8413_6 ( .COUTY1(na8413_4), .COUTY2(na8413_5), .POUTY1(na8413_7), .CINX(na8403_3), .CINY1(na8412_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na8412_7), .PINY2(1'b0), .OUT1(na8413_1), .OUT2(1'b0), .COMP_OUT(na8413_3_i) );
// C_MULTFa//O_O2//      x131y107     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a8414_1 ( .COUTY1(na8414_4), .COUTY2(na8414_5), .POUTY1(na8414_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1),
                      .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na8404_3), .CINY1(na8413_4), .CINY2(na8413_5),
                      .PINX(1'b0), .PINY1(na8413_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x131y108     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a8415_1 ( .OUT(na8415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na8414_4), .PINX(1'b0), .PINY1(na8414_7) );
C_O_0      #(.CPE_CFG ()) 
           _a8415_3 ( .COMP_OUT(na8415_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a8415_4 ( .OUT(na8415_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na8414_4), .PINX(1'b0), .PINY1(na8414_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a8415_6 ( .COUTY1(na8415_4), .COUTY2(na8415_5), .POUTY1(na8415_7), .POUTY2(na8415_8), .CINX(1'b0), .CINY1(na8414_4), .CINY2(na8414_5),
                      .PINX(1'b0), .PINY1(na8414_7), .PINY2(1'b0), .OUT1(na8415_1), .OUT2(na8415_2), .COMP_OUT(na8415_3_i) );
// C_MULT///MULT/      x131y109     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8416_1 ( .OUT1(na8416_1), .OUT2(na8416_2), .COUTY1(na8416_4), .COUTY2(na8416_5), .POUTY1(na8416_7), .POUTY2(na8416_8), .IN1(na8384_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na8384_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8383_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na8406_3), .CINY1(na8415_4), .CINY2(na8415_5), .PINX(na8406_6), .PINY1(na8415_7), .PINY2(na8415_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x131y110     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8417_1 ( .OUT1(na8417_1), .COUTY1(na8417_4), .COUTY2(na8417_5), .POUTY1(na8417_7), .POUTY2(na8417_8), .IN1(~na8385_2), .IN2(1'b1),
                      .IN3(1'b1), .IN4(1'b1), .IN5(~na8385_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8384_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0),
                      .CINX(na8407_3), .CINY1(na8416_4), .CINY2(na8416_5), .PINX(na8407_6), .PINY1(na8416_7), .PINY2(na8416_8), .RAM_I1(1'b0),
                      .RAM_I2(1'b0) );
// C_MULT///MULT/      x131y111     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8418_1 ( .COUTY1(na8418_4), .COUTY2(na8418_5), .POUTY1(na8418_7), .POUTY2(na8418_8), .IN1(na8386_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na8386_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8385_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na8408_3),
                      .CINY1(na8417_4), .CINY2(na8417_5), .PINX(na8408_6), .PINY1(na8417_7), .PINY2(na8417_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x131y112     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8419_1 ( .COUTY1(na8419_4), .COUTY2(na8419_5), .POUTY1(na8419_7), .POUTY2(na8419_8), .IN1(~na8387_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na8387_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8386_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na8409_3),
                      .CINY1(na8418_4), .CINY2(na8418_5), .PINX(na8409_6), .PINY1(na8418_7), .PINY2(na8418_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x131y113     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a8420_1 ( .COUTY1(na8420_4), .COUTY2(na8420_5), .POUTY1(na8420_7), .POUTY2(na8420_8), .IN1(na8388_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na8388_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na8387_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na8410_3),
                      .CINY1(na8419_4), .CINY2(na8419_5), .PINX(na8410_6), .PINY1(na8419_7), .PINY2(na8419_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x131y114     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a8421_1 ( .COUTY1(na8421_4), .COUTY2(na8421_5), .POUTY1(na8421_7), .POUTY2(na8421_8), .IN1(~na8389_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na8389_1), .IN6(1'b1), .IN7(1'b1), .IN8(na8388_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na8411_3),
                      .CINY1(na8420_4), .CINY2(na8420_5), .PINX(na8411_6), .PINY1(na8420_7), .PINY2(na8420_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x131y115     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a8422_3 ( .COMP_OUT(na8422_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a8422_4 ( .OUT(na8422_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na8421_4), .PINX(1'b0), .PINY1(na8421_7) );
// C_///AND/      x69y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8423_4 ( .OUT(na8423_2), .IN1(1'b1), .IN2(na1880_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8423_6 ( .RAM_O2(na8423_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8423_2), .COMP_OUT(1'b0) );
// C_///AND/      x85y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8424_4 ( .OUT(na8424_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1061_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8424_6 ( .RAM_O2(na8424_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8424_2), .COMP_OUT(1'b0) );
// C_///AND/      x86y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8425_4 ( .OUT(na8425_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1061_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8425_6 ( .RAM_O2(na8425_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8425_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y83     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8426_4 ( .OUT(na8426_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2818_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8426_6 ( .RAM_O2(na8426_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8426_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y84     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8427_4 ( .OUT(na8427_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2818_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8427_6 ( .RAM_O2(na8427_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8427_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y77     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8428_4 ( .OUT(na8428_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2805_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8428_6 ( .RAM_O2(na8428_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8428_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y78     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8429_4 ( .OUT(na8429_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2805_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8429_6 ( .RAM_O2(na8429_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8429_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y79     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8430_4 ( .OUT(na8430_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2811_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8430_6 ( .RAM_O2(na8430_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8430_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y80     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8431_4 ( .OUT(na8431_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2811_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8431_6 ( .RAM_O2(na8431_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8431_2), .COMP_OUT(1'b0) );
// C_///AND/      x123y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8432_4 ( .OUT(na8432_2), .IN1(1'b1), .IN2(1'b1), .IN3(na4930_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8432_6 ( .RAM_O2(na8432_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8432_2), .COMP_OUT(1'b0) );
// C_///AND/      x121y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8433_4 ( .OUT(na8433_2), .IN1(na4926_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8433_6 ( .RAM_O2(na8433_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8433_2), .COMP_OUT(1'b0) );
// C_///AND/      x109y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8434_4 ( .OUT(na8434_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2986_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8434_6 ( .RAM_O2(na8434_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8434_2), .COMP_OUT(1'b0) );
// C_///AND/      x113y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8435_4 ( .OUT(na8435_2), .IN1(1'b1), .IN2(na4936_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8435_6 ( .RAM_O2(na8435_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8435_2), .COMP_OUT(1'b0) );
// C_///AND/      x114y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8436_4 ( .OUT(na8436_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8436_6 ( .RAM_O2(na8436_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8436_2), .COMP_OUT(1'b0) );
// C_///AND/      x125y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8437_4 ( .OUT(na8437_2), .IN1(1'b1), .IN2(na4860_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8437_6 ( .RAM_O2(na8437_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8437_2), .COMP_OUT(1'b0) );
// C_///AND/      x126y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8438_4 ( .OUT(na8438_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8438_6 ( .RAM_O2(na8438_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8438_2), .COMP_OUT(1'b0) );
// C_///AND/      x117y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8439_4 ( .OUT(na8439_2), .IN1(na4864_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8439_6 ( .RAM_O2(na8439_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8439_2), .COMP_OUT(1'b0) );
// C_///AND/      x118y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8440_4 ( .OUT(na8440_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8440_6 ( .RAM_O2(na8440_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8440_2), .COMP_OUT(1'b0) );
// C_///AND/      x119y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8441_4 ( .OUT(na8441_2), .IN1(1'b1), .IN2(na4868_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8441_6 ( .RAM_O2(na8441_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8441_2), .COMP_OUT(1'b0) );
// C_///AND/      x120y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8442_4 ( .OUT(na8442_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8442_6 ( .RAM_O2(na8442_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8442_2), .COMP_OUT(1'b0) );
// C_///AND/      x103y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8443_4 ( .OUT(na8443_2), .IN1(1'b1), .IN2(na4872_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8443_6 ( .RAM_O2(na8443_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8443_2), .COMP_OUT(1'b0) );
// C_///AND/      x104y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8444_4 ( .OUT(na8444_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8444_6 ( .RAM_O2(na8444_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8444_2), .COMP_OUT(1'b0) );
// C_///AND/      x105y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8445_4 ( .OUT(na8445_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4876_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8445_6 ( .RAM_O2(na8445_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8445_2), .COMP_OUT(1'b0) );
// C_///AND/      x106y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8446_4 ( .OUT(na8446_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8446_6 ( .RAM_O2(na8446_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8446_2), .COMP_OUT(1'b0) );
// C_///AND/      x127y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8447_4 ( .OUT(na8447_2), .IN1(1'b1), .IN2(1'b1), .IN3(na4882_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8447_6 ( .RAM_O2(na8447_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8447_2), .COMP_OUT(1'b0) );
// C_///AND/      x128y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8448_4 ( .OUT(na8448_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8448_6 ( .RAM_O2(na8448_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8448_2), .COMP_OUT(1'b0) );
// C_///AND/      x135y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8449_4 ( .OUT(na8449_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4886_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8449_6 ( .RAM_O2(na8449_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8449_2), .COMP_OUT(1'b0) );
// C_///AND/      x136y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8450_4 ( .OUT(na8450_2), .IN1(na4933_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8450_6 ( .RAM_O2(na8450_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8450_2), .COMP_OUT(1'b0) );
// C_///AND/      x101y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8451_4 ( .OUT(na8451_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2789_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8451_6 ( .RAM_O2(na8451_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8451_2), .COMP_OUT(1'b0) );
// C_///AND/      x111y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8452_4 ( .OUT(na8452_2), .IN1(na4893_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8452_6 ( .RAM_O2(na8452_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8452_2), .COMP_OUT(1'b0) );
// C_///AND/      x112y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8453_4 ( .OUT(na8453_2), .IN1(na4890_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8453_6 ( .RAM_O2(na8453_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8453_2), .COMP_OUT(1'b0) );
// C_///AND/      x77y1     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8454_4 ( .OUT(na8454_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8454_6 ( .RAM_O2(na8454_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8454_2), .COMP_OUT(1'b0) );
// C_///AND/      x78y1     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8455_4 ( .OUT(na8455_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na2699_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8455_6 ( .RAM_O2(na8455_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8455_2), .COMP_OUT(1'b0) );
// C_///AND/      x79y1     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8456_4 ( .OUT(na8456_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8456_6 ( .RAM_O2(na8456_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8456_2), .COMP_OUT(1'b0) );
// C_///AND/      x80y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8457_4 ( .OUT(na8457_2), .IN1(1'b1), .IN2(1'b1), .IN3(na5_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8457_6 ( .RAM_O2(na8457_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8457_2), .COMP_OUT(1'b0) );
// C_///AND/      x85y1     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8458_4 ( .OUT(na8458_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8458_6 ( .RAM_O2(na8458_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8458_2), .COMP_OUT(1'b0) );
// C_///AND/      x86y1     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8459_4 ( .OUT(na8459_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na2698_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8459_6 ( .RAM_O2(na8459_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8459_2), .COMP_OUT(1'b0) );
// C_///AND/      x87y1     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8460_4 ( .OUT(na8460_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8460_6 ( .RAM_O2(na8460_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8460_2), .COMP_OUT(1'b0) );
// C_///AND/      x88y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8461_4 ( .OUT(na8461_2), .IN1(1'b1), .IN2(na6_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8461_6 ( .RAM_O2(na8461_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8461_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y39     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8462_4 ( .OUT(na8462_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1065_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8462_6 ( .RAM_O2(na8462_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8462_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y40     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8463_4 ( .OUT(na8463_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1065_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8463_6 ( .RAM_O2(na8463_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8463_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8464_4 ( .OUT(na8464_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2687_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8464_6 ( .RAM_O2(na8464_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8464_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y38     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8465_4 ( .OUT(na8465_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2687_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8465_6 ( .RAM_O2(na8465_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8465_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y47     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8466_4 ( .OUT(na8466_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1359_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8466_6 ( .RAM_O2(na8466_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8466_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y48     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8467_4 ( .OUT(na8467_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1359_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8467_6 ( .RAM_O2(na8467_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8467_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y45     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8468_4 ( .OUT(na8468_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1355_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8468_6 ( .RAM_O2(na8468_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8468_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y46     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8469_4 ( .OUT(na8469_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1355_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8469_6 ( .RAM_O2(na8469_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8469_2), .COMP_OUT(1'b0) );
// C_///AND/      x79y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8470_4 ( .OUT(na8470_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2681_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8470_6 ( .RAM_O2(na8470_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8470_2), .COMP_OUT(1'b0) );
// C_///AND/      x80y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8471_4 ( .OUT(na8471_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2681_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8471_6 ( .RAM_O2(na8471_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8471_2), .COMP_OUT(1'b0) );
// C_///AND/      x59y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8472_4 ( .OUT(na8472_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1314_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8472_6 ( .RAM_O2(na8472_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8472_2), .COMP_OUT(1'b0) );
// C_///AND/      x60y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8473_4 ( .OUT(na8473_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1314_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8473_6 ( .RAM_O2(na8473_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8473_2), .COMP_OUT(1'b0) );
// C_///AND/      x57y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8474_4 ( .OUT(na8474_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2677_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8474_6 ( .RAM_O2(na8474_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8474_2), .COMP_OUT(1'b0) );
// C_///AND/      x58y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8475_4 ( .OUT(na8475_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2677_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8475_6 ( .RAM_O2(na8475_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8475_2), .COMP_OUT(1'b0) );
// C_///AND/      x61y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8476_4 ( .OUT(na8476_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1337_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8476_6 ( .RAM_O2(na8476_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8476_2), .COMP_OUT(1'b0) );
// C_///AND/      x62y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8477_4 ( .OUT(na8477_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1337_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8477_6 ( .RAM_O2(na8477_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8477_2), .COMP_OUT(1'b0) );
// C_///AND/      x65y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8478_4 ( .OUT(na8478_2), .IN1(1'b1), .IN2(1'b1), .IN3(na913_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8478_6 ( .RAM_O2(na8478_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8478_2), .COMP_OUT(1'b0) );
// C_///AND/      x66y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8479_4 ( .OUT(na8479_2), .IN1(1'b1), .IN2(1'b1), .IN3(na913_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8479_6 ( .RAM_O2(na8479_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8479_2), .COMP_OUT(1'b0) );
// C_///AND/      x67y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8480_4 ( .OUT(na8480_2), .IN1(1'b1), .IN2(1'b1), .IN3(na925_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8480_6 ( .RAM_O2(na8480_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8480_2), .COMP_OUT(1'b0) );
// C_///AND/      x68y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8481_4 ( .OUT(na8481_2), .IN1(1'b1), .IN2(1'b1), .IN3(na925_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8481_6 ( .RAM_O2(na8481_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8481_2), .COMP_OUT(1'b0) );
// C_///AND/      x69y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8482_4 ( .OUT(na8482_2), .IN1(1'b1), .IN2(na927_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8482_6 ( .RAM_O2(na8482_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8482_2), .COMP_OUT(1'b0) );
// C_///AND/      x39y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8483_4 ( .OUT(na8483_2), .IN1(1'b1), .IN2(na2749_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8483_6 ( .RAM_O2(na8483_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8483_2), .COMP_OUT(1'b0) );
// C_///AND/      x37y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8484_4 ( .OUT(na8484_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2830_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8484_6 ( .RAM_O2(na8484_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8484_2), .COMP_OUT(1'b0) );
// C_///AND/      x35y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8485_4 ( .OUT(na8485_2), .IN1(1'b1), .IN2(na6090_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8485_6 ( .RAM_O2(na8485_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8485_2), .COMP_OUT(1'b0) );
// C_///AND/      x87y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8486_4 ( .OUT(na8486_2), .IN1(1'b1), .IN2(na2722_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8486_6 ( .RAM_O2(na8486_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8486_2), .COMP_OUT(1'b0) );
// C_///AND/      x75y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8487_4 ( .OUT(na8487_2), .IN1(1'b1), .IN2(1'b1), .IN3(na930_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8487_6 ( .RAM_O2(na8487_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8487_2), .COMP_OUT(1'b0) );
// C_///AND/      x73y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8488_4 ( .OUT(na8488_2), .IN1(na6004_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8488_6 ( .RAM_O2(na8488_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8488_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y25     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8489_4 ( .OUT(na8489_2), .IN1(na3588_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8489_6 ( .RAM_O2(na8489_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8489_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y53     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8490_4 ( .OUT(na8490_2), .IN1(1'b1), .IN2(1'b1), .IN3(na3548_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8490_6 ( .RAM_O2(na8490_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8490_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y85     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8491_4 ( .OUT(na8491_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1409_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8491_6 ( .RAM_O2(na8491_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8491_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y27     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8492_4 ( .OUT(na8492_2), .IN1(1'b1), .IN2(1'b1), .IN3(na945_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8492_6 ( .RAM_O2(na8492_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8492_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y31     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8493_4 ( .OUT(na8493_2), .IN1(na948_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8493_6 ( .RAM_O2(na8493_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8493_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y25     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8494_4 ( .OUT(na8494_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na949_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8494_6 ( .RAM_O2(na8494_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8494_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y29     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8495_4 ( .OUT(na8495_2), .IN1(1'b1), .IN2(na958_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8495_6 ( .RAM_O2(na8495_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8495_2), .COMP_OUT(1'b0) );
// C_///AND/      x71y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8496_4 ( .OUT(na8496_2), .IN1(1'b1), .IN2(na942_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8496_6 ( .RAM_O2(na8496_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8496_2), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y64     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8497_4 ( .OUT(na8497_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8497_5 ( .OUT(na8497_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8497_6 ( .RAM_O2(na8497_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8497_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y64     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8498_1 ( .OUT(na8498_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8498_2 ( .OUT(na8498_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8498_6 ( .RAM_O1(na8498_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8498_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y63     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8499_4 ( .OUT(na8499_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8499_5 ( .OUT(na8499_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8499_6 ( .RAM_O2(na8499_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8499_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y63     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8500_1 ( .OUT(na8500_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8500_2 ( .OUT(na8500_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8500_6 ( .RAM_O1(na8500_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8500_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y62     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8501_4 ( .OUT(na8501_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8501_5 ( .OUT(na8501_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8501_6 ( .RAM_O2(na8501_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8501_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y62     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8502_1 ( .OUT(na8502_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8502_2 ( .OUT(na8502_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8502_6 ( .RAM_O1(na8502_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8502_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y61     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8503_4 ( .OUT(na8503_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8503_5 ( .OUT(na8503_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8503_6 ( .RAM_O2(na8503_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8503_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y61     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8504_1 ( .OUT(na8504_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8504_2 ( .OUT(na8504_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8504_6 ( .RAM_O1(na8504_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8504_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y60     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8505_4 ( .OUT(na8505_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8505_5 ( .OUT(na8505_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8505_6 ( .RAM_O2(na8505_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8505_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y60     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8506_1 ( .OUT(na8506_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8506_2 ( .OUT(na8506_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8506_6 ( .RAM_O1(na8506_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8506_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y59     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8507_4 ( .OUT(na8507_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8507_5 ( .OUT(na8507_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8507_6 ( .RAM_O2(na8507_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8507_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y59     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8508_1 ( .OUT(na8508_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8508_2 ( .OUT(na8508_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8508_6 ( .RAM_O1(na8508_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8508_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y58     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8509_4 ( .OUT(na8509_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8509_5 ( .OUT(na8509_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8509_6 ( .RAM_O2(na8509_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8509_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y58     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8510_1 ( .OUT(na8510_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8510_2 ( .OUT(na8510_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8510_6 ( .RAM_O1(na8510_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8510_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y57     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8511_4 ( .OUT(na8511_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8511_5 ( .OUT(na8511_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8511_6 ( .RAM_O2(na8511_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8511_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y57     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8512_1 ( .OUT(na8512_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8512_2 ( .OUT(na8512_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8512_6 ( .RAM_O1(na8512_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8512_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y52     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8513_4 ( .OUT(na8513_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8513_5 ( .OUT(na8513_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8513_6 ( .RAM_O2(na8513_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8513_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y52     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8514_1 ( .OUT(na8514_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8514_2 ( .OUT(na8514_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8514_6 ( .RAM_O1(na8514_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8514_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y51     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8515_4 ( .OUT(na8515_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8515_5 ( .OUT(na8515_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8515_6 ( .RAM_O2(na8515_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8515_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y51     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8516_1 ( .OUT(na8516_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8516_2 ( .OUT(na8516_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8516_6 ( .RAM_O1(na8516_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8516_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y50     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8517_4 ( .OUT(na8517_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8517_5 ( .OUT(na8517_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8517_6 ( .RAM_O2(na8517_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8517_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y50     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8518_1 ( .OUT(na8518_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8518_2 ( .OUT(na8518_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8518_6 ( .RAM_O1(na8518_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8518_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y49     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8519_4 ( .OUT(na8519_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8519_5 ( .OUT(na8519_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8519_6 ( .RAM_O2(na8519_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8519_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y49     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8520_1 ( .OUT(na8520_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8520_2 ( .OUT(na8520_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6650_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8520_6 ( .RAM_O1(na8520_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8520_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y64     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8521_4 ( .OUT(na8521_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2866_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8521_6 ( .RAM_O2(na8521_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8521_2), .COMP_OUT(1'b0) );
// C_AND////      x29y64     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8522_1 ( .OUT(na8522_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2866_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8522_6 ( .RAM_O1(na8522_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8522_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y63     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8523_4 ( .OUT(na8523_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2866_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8523_6 ( .RAM_O2(na8523_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8523_2), .COMP_OUT(1'b0) );
// C_AND////      x29y63     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8524_1 ( .OUT(na8524_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2866_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8524_6 ( .RAM_O1(na8524_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8524_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y64     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8525_4 ( .OUT(na8525_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2866_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8525_6 ( .RAM_O2(na8525_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8525_2), .COMP_OUT(1'b0) );
// C_AND////      x31y64     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8526_1 ( .OUT(na8526_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2866_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8526_6 ( .RAM_O1(na8526_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8526_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y63     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8527_4 ( .OUT(na8527_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2866_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8527_6 ( .RAM_O2(na8527_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8527_2), .COMP_OUT(1'b0) );
// C_AND////      x31y63     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8528_1 ( .OUT(na8528_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2866_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8528_6 ( .RAM_O1(na8528_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8528_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y62     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8529_4 ( .OUT(na8529_2), .IN1(1'b1), .IN2(na2865_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8529_6 ( .RAM_O2(na8529_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8529_2), .COMP_OUT(1'b0) );
// C_AND////      x31y62     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8530_1 ( .OUT(na8530_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2865_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8530_6 ( .RAM_O1(na8530_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8530_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y61     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8531_4 ( .OUT(na8531_2), .IN1(1'b1), .IN2(na2865_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8531_6 ( .RAM_O2(na8531_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8531_2), .COMP_OUT(1'b0) );
// C_AND////      x31y61     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8532_1 ( .OUT(na8532_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2865_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8532_6 ( .RAM_O1(na8532_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8532_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y60     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8533_4 ( .OUT(na8533_2), .IN1(1'b1), .IN2(na2865_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8533_6 ( .RAM_O2(na8533_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8533_2), .COMP_OUT(1'b0) );
// C_AND////      x31y60     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8534_1 ( .OUT(na8534_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2865_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8534_6 ( .RAM_O1(na8534_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8534_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y59     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8535_4 ( .OUT(na8535_2), .IN1(1'b1), .IN2(na2865_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8535_6 ( .RAM_O2(na8535_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8535_2), .COMP_OUT(1'b0) );
// C_AND////      x31y59     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8536_1 ( .OUT(na8536_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2865_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8536_6 ( .RAM_O1(na8536_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8536_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y58     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8537_4 ( .OUT(na8537_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2863_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8537_6 ( .RAM_O2(na8537_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8537_2), .COMP_OUT(1'b0) );
// C_AND////      x31y58     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8538_1 ( .OUT(na8538_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2863_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8538_6 ( .RAM_O1(na8538_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8538_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y57     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8539_4 ( .OUT(na8539_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2863_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8539_6 ( .RAM_O2(na8539_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8539_2), .COMP_OUT(1'b0) );
// C_AND////      x31y57     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8540_1 ( .OUT(na8540_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2863_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8540_6 ( .RAM_O1(na8540_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8540_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x35y73     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8541_1 ( .OUT(na8541_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8541_6 ( .RAM_O1(na8541_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8541_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x35y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8542_1 ( .OUT(na8542_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8542_6 ( .RAM_O1(na8542_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8542_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y73     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8543_4 ( .OUT(na8543_2), .IN1(1'b1), .IN2(na3231_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8543_6 ( .RAM_O2(na8543_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8543_2), .COMP_OUT(1'b0) );
// C_///AND/      x27y65     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8544_4 ( .OUT(na8544_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3233_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8544_6 ( .RAM_O2(na8544_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8544_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y72     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8545_4 ( .OUT(na8545_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8545_6 ( .RAM_O2(na8545_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8545_2), .COMP_OUT(1'b0) );
// C_AND////      x28y72     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8546_1 ( .OUT(na8546_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8546_6 ( .RAM_O1(na8546_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8546_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y71     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8547_4 ( .OUT(na8547_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8547_6 ( .RAM_O2(na8547_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8547_2), .COMP_OUT(1'b0) );
// C_AND////      x28y71     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8548_1 ( .OUT(na8548_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8548_6 ( .RAM_O1(na8548_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8548_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y70     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8549_4 ( .OUT(na8549_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8549_6 ( .RAM_O2(na8549_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8549_2), .COMP_OUT(1'b0) );
// C_AND////      x28y70     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8550_1 ( .OUT(na8550_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8550_6 ( .RAM_O1(na8550_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8550_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y69     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8551_4 ( .OUT(na8551_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8551_6 ( .RAM_O2(na8551_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8551_2), .COMP_OUT(1'b0) );
// C_AND////      x28y69     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8552_1 ( .OUT(na8552_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8552_6 ( .RAM_O1(na8552_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8552_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y68     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8553_4 ( .OUT(na8553_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8553_6 ( .RAM_O2(na8553_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8553_2), .COMP_OUT(1'b0) );
// C_AND////      x28y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8554_1 ( .OUT(na8554_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8554_6 ( .RAM_O1(na8554_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8554_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y67     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8555_4 ( .OUT(na8555_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8555_6 ( .RAM_O2(na8555_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8555_2), .COMP_OUT(1'b0) );
// C_AND////      x28y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8556_1 ( .OUT(na8556_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8556_6 ( .RAM_O1(na8556_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8556_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8557_4 ( .OUT(na8557_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8557_6 ( .RAM_O2(na8557_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8557_2), .COMP_OUT(1'b0) );
// C_AND////      x28y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8558_1 ( .OUT(na8558_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8558_6 ( .RAM_O1(na8558_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8558_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8559_4 ( .OUT(na8559_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8559_6 ( .RAM_O2(na8559_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8559_2), .COMP_OUT(1'b0) );
// C_AND////      x28y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8560_1 ( .OUT(na8560_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8560_6 ( .RAM_O1(na8560_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8560_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y80     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8561_4 ( .OUT(na8561_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8561_6 ( .RAM_O2(na8561_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8561_2), .COMP_OUT(1'b0) );
// C_AND////      x28y80     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8562_1 ( .OUT(na8562_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8562_6 ( .RAM_O1(na8562_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8562_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y79     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8563_4 ( .OUT(na8563_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8563_6 ( .RAM_O2(na8563_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8563_2), .COMP_OUT(1'b0) );
// C_AND////      x28y79     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8564_1 ( .OUT(na8564_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8564_6 ( .RAM_O1(na8564_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8564_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y78     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8565_4 ( .OUT(na8565_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8565_6 ( .RAM_O2(na8565_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8565_2), .COMP_OUT(1'b0) );
// C_AND////      x28y78     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8566_1 ( .OUT(na8566_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8566_6 ( .RAM_O1(na8566_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8566_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y77     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8567_4 ( .OUT(na8567_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8567_6 ( .RAM_O2(na8567_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8567_2), .COMP_OUT(1'b0) );
// C_AND////      x28y77     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8568_1 ( .OUT(na8568_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8568_6 ( .RAM_O1(na8568_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8568_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y76     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8569_4 ( .OUT(na8569_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8569_6 ( .RAM_O2(na8569_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8569_2), .COMP_OUT(1'b0) );
// C_AND////      x28y76     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8570_1 ( .OUT(na8570_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8570_6 ( .RAM_O1(na8570_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8570_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y75     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8571_4 ( .OUT(na8571_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8571_6 ( .RAM_O2(na8571_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8571_2), .COMP_OUT(1'b0) );
// C_AND////      x28y75     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8572_1 ( .OUT(na8572_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8572_6 ( .RAM_O1(na8572_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8572_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y74     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8573_4 ( .OUT(na8573_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8573_6 ( .RAM_O2(na8573_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8573_2), .COMP_OUT(1'b0) );
// C_AND////      x28y74     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8574_1 ( .OUT(na8574_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8574_6 ( .RAM_O1(na8574_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8574_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y73     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8575_4 ( .OUT(na8575_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8575_6 ( .RAM_O2(na8575_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8575_2), .COMP_OUT(1'b0) );
// C_AND////      x28y73     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8576_1 ( .OUT(na8576_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8576_6 ( .RAM_O1(na8576_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8576_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x37y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8577_1 ( .OUT(na8577_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8577_6 ( .RAM_O1(na8577_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8577_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x37y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8578_1 ( .OUT(na8578_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8578_6 ( .RAM_O1(na8578_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8578_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8579_4 ( .OUT(na8579_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8579_6 ( .RAM_O2(na8579_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8579_2), .COMP_OUT(1'b0) );
// C_AND////      x37y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8580_1 ( .OUT(na8580_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8580_6 ( .RAM_O1(na8580_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8580_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8581_4 ( .OUT(na8581_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8581_6 ( .RAM_O2(na8581_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8581_2), .COMP_OUT(1'b0) );
// C_AND////      x37y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8582_1 ( .OUT(na8582_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8582_6 ( .RAM_O1(na8582_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8582_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x37y76     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8583_1 ( .OUT(na8583_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8583_6 ( .RAM_O1(na8583_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8583_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x37y75     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8584_1 ( .OUT(na8584_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8584_6 ( .RAM_O1(na8584_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8584_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y74     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8585_4 ( .OUT(na8585_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8585_6 ( .RAM_O2(na8585_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8585_2), .COMP_OUT(1'b0) );
// C_AND////      x37y74     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8586_1 ( .OUT(na8586_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8586_6 ( .RAM_O1(na8586_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8586_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y73     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8587_4 ( .OUT(na8587_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8587_6 ( .RAM_O2(na8587_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8587_2), .COMP_OUT(1'b0) );
// C_AND////      x37y73     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8588_1 ( .OUT(na8588_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8588_6 ( .RAM_O1(na8588_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8588_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x30y80     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8589_4 ( .OUT(na8589_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8589_5 ( .OUT(na8589_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8589_6 ( .RAM_O2(na8589_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8589_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x30y80     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8590_1 ( .OUT(na8590_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8590_2 ( .OUT(na8590_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8590_6 ( .RAM_O1(na8590_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8590_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x30y79     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8591_4 ( .OUT(na8591_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8591_5 ( .OUT(na8591_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8591_6 ( .RAM_O2(na8591_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8591_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x30y79     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8592_1 ( .OUT(na8592_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8592_2 ( .OUT(na8592_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8592_6 ( .RAM_O1(na8592_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8592_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y80     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8593_4 ( .OUT(na8593_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8593_5 ( .OUT(na8593_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8593_6 ( .RAM_O2(na8593_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8593_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y80     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8594_1 ( .OUT(na8594_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8594_2 ( .OUT(na8594_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8594_6 ( .RAM_O1(na8594_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8594_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y79     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8595_4 ( .OUT(na8595_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8595_5 ( .OUT(na8595_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8595_6 ( .RAM_O2(na8595_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8595_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y79     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8596_1 ( .OUT(na8596_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8596_2 ( .OUT(na8596_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8596_6 ( .RAM_O1(na8596_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8596_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y78     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8597_4 ( .OUT(na8597_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8597_5 ( .OUT(na8597_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8597_6 ( .RAM_O2(na8597_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8597_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y78     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8598_1 ( .OUT(na8598_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8598_2 ( .OUT(na8598_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8598_6 ( .RAM_O1(na8598_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8598_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y77     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8599_4 ( .OUT(na8599_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8599_5 ( .OUT(na8599_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8599_6 ( .RAM_O2(na8599_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8599_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y77     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8600_1 ( .OUT(na8600_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8600_2 ( .OUT(na8600_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8600_6 ( .RAM_O1(na8600_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8600_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y76     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8601_4 ( .OUT(na8601_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8601_5 ( .OUT(na8601_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8601_6 ( .RAM_O2(na8601_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8601_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y76     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8602_1 ( .OUT(na8602_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8602_2 ( .OUT(na8602_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8602_6 ( .RAM_O1(na8602_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8602_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y75     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8603_4 ( .OUT(na8603_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8603_5 ( .OUT(na8603_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8603_6 ( .RAM_O2(na8603_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8603_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y75     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8604_1 ( .OUT(na8604_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8604_2 ( .OUT(na8604_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8604_6 ( .RAM_O1(na8604_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8604_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y74     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8605_4 ( .OUT(na8605_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8605_5 ( .OUT(na8605_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8605_6 ( .RAM_O2(na8605_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8605_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y74     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8606_1 ( .OUT(na8606_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8606_2 ( .OUT(na8606_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8606_6 ( .RAM_O1(na8606_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8606_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y73     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8607_4 ( .OUT(na8607_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8607_5 ( .OUT(na8607_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8607_6 ( .RAM_O2(na8607_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8607_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y73     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8608_1 ( .OUT(na8608_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8608_2 ( .OUT(na8608_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8608_6 ( .RAM_O1(na8608_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8608_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x30y72     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8609_4 ( .OUT(na8609_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8609_5 ( .OUT(na8609_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8609_6 ( .RAM_O2(na8609_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8609_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x30y72     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8610_1 ( .OUT(na8610_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8610_2 ( .OUT(na8610_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8610_6 ( .RAM_O1(na8610_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8610_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x30y71     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8611_4 ( .OUT(na8611_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8611_5 ( .OUT(na8611_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8611_6 ( .RAM_O2(na8611_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8611_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x30y71     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8612_1 ( .OUT(na8612_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8612_2 ( .OUT(na8612_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8612_6 ( .RAM_O1(na8612_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8612_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y72     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8613_4 ( .OUT(na8613_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8613_5 ( .OUT(na8613_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8613_6 ( .RAM_O2(na8613_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8613_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y72     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8614_1 ( .OUT(na8614_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8614_2 ( .OUT(na8614_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8614_6 ( .RAM_O1(na8614_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8614_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y71     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8615_4 ( .OUT(na8615_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8615_5 ( .OUT(na8615_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8615_6 ( .RAM_O2(na8615_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8615_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y71     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8616_1 ( .OUT(na8616_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8616_2 ( .OUT(na8616_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8616_6 ( .RAM_O1(na8616_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8616_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y70     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8617_4 ( .OUT(na8617_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8617_5 ( .OUT(na8617_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8617_6 ( .RAM_O2(na8617_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8617_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y70     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8618_1 ( .OUT(na8618_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8618_2 ( .OUT(na8618_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8618_6 ( .RAM_O1(na8618_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8618_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y69     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8619_4 ( .OUT(na8619_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8619_5 ( .OUT(na8619_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8619_6 ( .RAM_O2(na8619_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8619_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y69     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8620_1 ( .OUT(na8620_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8620_2 ( .OUT(na8620_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8620_6 ( .RAM_O1(na8620_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8620_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y68     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8621_4 ( .OUT(na8621_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8621_5 ( .OUT(na8621_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8621_6 ( .RAM_O2(na8621_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8621_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y68     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8622_1 ( .OUT(na8622_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8622_2 ( .OUT(na8622_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8622_6 ( .RAM_O1(na8622_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8622_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y67     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8623_4 ( .OUT(na8623_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8623_5 ( .OUT(na8623_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8623_6 ( .RAM_O2(na8623_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8623_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y67     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8624_1 ( .OUT(na8624_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8624_2 ( .OUT(na8624_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8624_6 ( .RAM_O1(na8624_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8624_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y66     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8625_4 ( .OUT(na8625_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8625_5 ( .OUT(na8625_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8625_6 ( .RAM_O2(na8625_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8625_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y66     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8626_1 ( .OUT(na8626_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8626_2 ( .OUT(na8626_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8626_6 ( .RAM_O1(na8626_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8626_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y65     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8627_4 ( .OUT(na8627_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8627_5 ( .OUT(na8627_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8627_6 ( .RAM_O2(na8627_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8627_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y65     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8628_1 ( .OUT(na8628_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8628_2 ( .OUT(na8628_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6651_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8628_6 ( .RAM_O1(na8628_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8628_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y80     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8629_4 ( .OUT(na8629_2), .IN1(na2860_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8629_6 ( .RAM_O2(na8629_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8629_2), .COMP_OUT(1'b0) );
// C_AND////      x29y80     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8630_1 ( .OUT(na8630_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2860_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8630_6 ( .RAM_O1(na8630_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8630_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y79     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8631_4 ( .OUT(na8631_2), .IN1(na2860_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8631_6 ( .RAM_O2(na8631_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8631_2), .COMP_OUT(1'b0) );
// C_AND////      x29y79     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8632_1 ( .OUT(na8632_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2860_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8632_6 ( .RAM_O1(na8632_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8632_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y80     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8633_4 ( .OUT(na8633_2), .IN1(na2860_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8633_6 ( .RAM_O2(na8633_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8633_2), .COMP_OUT(1'b0) );
// C_AND////      x31y80     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8634_1 ( .OUT(na8634_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2860_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8634_6 ( .RAM_O1(na8634_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8634_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y79     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8635_4 ( .OUT(na8635_2), .IN1(na2860_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8635_6 ( .RAM_O2(na8635_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8635_2), .COMP_OUT(1'b0) );
// C_AND////      x31y79     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8636_1 ( .OUT(na8636_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2860_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8636_6 ( .RAM_O1(na8636_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8636_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y78     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8637_4 ( .OUT(na8637_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2858_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8637_6 ( .RAM_O2(na8637_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8637_2), .COMP_OUT(1'b0) );
// C_AND////      x31y78     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8638_1 ( .OUT(na8638_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2858_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8638_6 ( .RAM_O1(na8638_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8638_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y77     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8639_4 ( .OUT(na8639_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2858_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8639_6 ( .RAM_O2(na8639_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8639_2), .COMP_OUT(1'b0) );
// C_AND////      x31y77     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8640_1 ( .OUT(na8640_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2858_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8640_6 ( .RAM_O1(na8640_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8640_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y76     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8641_4 ( .OUT(na8641_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2858_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8641_6 ( .RAM_O2(na8641_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8641_2), .COMP_OUT(1'b0) );
// C_AND////      x31y76     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8642_1 ( .OUT(na8642_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2858_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8642_6 ( .RAM_O1(na8642_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8642_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y75     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8643_4 ( .OUT(na8643_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2858_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8643_6 ( .RAM_O2(na8643_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8643_2), .COMP_OUT(1'b0) );
// C_AND////      x31y75     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8644_1 ( .OUT(na8644_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2858_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8644_6 ( .RAM_O1(na8644_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8644_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y74     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8645_4 ( .OUT(na8645_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2857_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8645_6 ( .RAM_O2(na8645_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8645_2), .COMP_OUT(1'b0) );
// C_AND////      x31y74     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8646_1 ( .OUT(na8646_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2857_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8646_6 ( .RAM_O1(na8646_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8646_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y73     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8647_4 ( .OUT(na8647_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2857_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8647_6 ( .RAM_O2(na8647_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8647_2), .COMP_OUT(1'b0) );
// C_AND////      x31y73     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8648_1 ( .OUT(na8648_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2857_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8648_6 ( .RAM_O1(na8648_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8648_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y72     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8649_4 ( .OUT(na8649_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2857_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8649_6 ( .RAM_O2(na8649_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8649_2), .COMP_OUT(1'b0) );
// C_AND////      x29y72     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8650_1 ( .OUT(na8650_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2857_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8650_6 ( .RAM_O1(na8650_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8650_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y71     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8651_4 ( .OUT(na8651_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2857_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8651_6 ( .RAM_O2(na8651_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8651_2), .COMP_OUT(1'b0) );
// C_AND////      x29y71     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8652_1 ( .OUT(na8652_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2857_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8652_6 ( .RAM_O1(na8652_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8652_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y72     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8653_4 ( .OUT(na8653_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2856_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8653_6 ( .RAM_O2(na8653_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8653_2), .COMP_OUT(1'b0) );
// C_AND////      x31y72     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8654_1 ( .OUT(na8654_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2856_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8654_6 ( .RAM_O1(na8654_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8654_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y71     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8655_4 ( .OUT(na8655_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2856_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8655_6 ( .RAM_O2(na8655_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8655_2), .COMP_OUT(1'b0) );
// C_AND////      x31y71     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8656_1 ( .OUT(na8656_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2856_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8656_6 ( .RAM_O1(na8656_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8656_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y70     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8657_4 ( .OUT(na8657_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2856_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8657_6 ( .RAM_O2(na8657_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8657_2), .COMP_OUT(1'b0) );
// C_AND////      x31y70     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8658_1 ( .OUT(na8658_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2856_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8658_6 ( .RAM_O1(na8658_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8658_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y69     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8659_4 ( .OUT(na8659_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2856_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8659_6 ( .RAM_O2(na8659_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8659_2), .COMP_OUT(1'b0) );
// C_AND////      x31y69     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8660_1 ( .OUT(na8660_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2856_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8660_6 ( .RAM_O1(na8660_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8660_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y68     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8661_4 ( .OUT(na8661_2), .IN1(na2855_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8661_6 ( .RAM_O2(na8661_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8661_2), .COMP_OUT(1'b0) );
// C_AND////      x31y68     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8662_1 ( .OUT(na8662_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2855_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8662_6 ( .RAM_O1(na8662_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8662_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y67     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8663_4 ( .OUT(na8663_2), .IN1(na2855_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8663_6 ( .RAM_O2(na8663_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8663_2), .COMP_OUT(1'b0) );
// C_AND////      x31y67     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8664_1 ( .OUT(na8664_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2855_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8664_6 ( .RAM_O1(na8664_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8664_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y66     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8665_4 ( .OUT(na8665_2), .IN1(na2855_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8665_6 ( .RAM_O2(na8665_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8665_2), .COMP_OUT(1'b0) );
// C_AND////      x31y66     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8666_1 ( .OUT(na8666_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2855_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8666_6 ( .RAM_O1(na8666_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8666_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y65     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8667_4 ( .OUT(na8667_2), .IN1(na2855_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8667_6 ( .RAM_O2(na8667_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8667_2), .COMP_OUT(1'b0) );
// C_AND////      x31y65     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8668_1 ( .OUT(na8668_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2855_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8668_6 ( .RAM_O1(na8668_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8668_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x67y25     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8669_1 ( .OUT(na8669_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8669_6 ( .RAM_O1(na8669_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8669_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x67y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8670_1 ( .OUT(na8670_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8670_6 ( .RAM_O1(na8670_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8670_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x59y25     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8671_4 ( .OUT(na8671_2), .IN1(1'b1), .IN2(na3303_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8671_6 ( .RAM_O2(na8671_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8671_2), .COMP_OUT(1'b0) );
// C_///AND/      x59y17     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8672_4 ( .OUT(na8672_2), .IN1(1'b1), .IN2(na3230_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8672_6 ( .RAM_O2(na8672_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8672_2), .COMP_OUT(1'b0) );
// C_///AND/      x60y24     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8673_4 ( .OUT(na8673_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8673_6 ( .RAM_O2(na8673_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8673_2), .COMP_OUT(1'b0) );
// C_AND////      x60y24     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8674_1 ( .OUT(na8674_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8674_6 ( .RAM_O1(na8674_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8674_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y23     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8675_4 ( .OUT(na8675_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8675_6 ( .RAM_O2(na8675_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8675_2), .COMP_OUT(1'b0) );
// C_AND////      x60y23     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8676_1 ( .OUT(na8676_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8676_6 ( .RAM_O1(na8676_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8676_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y22     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8677_4 ( .OUT(na8677_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8677_6 ( .RAM_O2(na8677_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8677_2), .COMP_OUT(1'b0) );
// C_AND////      x60y22     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8678_1 ( .OUT(na8678_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8678_6 ( .RAM_O1(na8678_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8678_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y21     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8679_4 ( .OUT(na8679_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8679_6 ( .RAM_O2(na8679_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8679_2), .COMP_OUT(1'b0) );
// C_AND////      x60y21     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8680_1 ( .OUT(na8680_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8680_6 ( .RAM_O1(na8680_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8680_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y20     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8681_4 ( .OUT(na8681_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8681_6 ( .RAM_O2(na8681_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8681_2), .COMP_OUT(1'b0) );
// C_AND////      x60y20     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8682_1 ( .OUT(na8682_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8682_6 ( .RAM_O1(na8682_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8682_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y19     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8683_4 ( .OUT(na8683_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8683_6 ( .RAM_O2(na8683_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8683_2), .COMP_OUT(1'b0) );
// C_AND////      x60y19     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8684_1 ( .OUT(na8684_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8684_6 ( .RAM_O1(na8684_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8684_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8685_4 ( .OUT(na8685_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8685_6 ( .RAM_O2(na8685_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8685_2), .COMP_OUT(1'b0) );
// C_AND////      x60y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8686_1 ( .OUT(na8686_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8686_6 ( .RAM_O1(na8686_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8686_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8687_4 ( .OUT(na8687_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8687_6 ( .RAM_O2(na8687_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8687_2), .COMP_OUT(1'b0) );
// C_AND////      x60y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8688_1 ( .OUT(na8688_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8688_6 ( .RAM_O1(na8688_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8688_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y32     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8689_4 ( .OUT(na8689_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8689_6 ( .RAM_O2(na8689_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8689_2), .COMP_OUT(1'b0) );
// C_AND////      x60y32     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8690_1 ( .OUT(na8690_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8690_6 ( .RAM_O1(na8690_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8690_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y31     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8691_4 ( .OUT(na8691_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8691_6 ( .RAM_O2(na8691_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8691_2), .COMP_OUT(1'b0) );
// C_AND////      x60y31     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8692_1 ( .OUT(na8692_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8692_6 ( .RAM_O1(na8692_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8692_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y30     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8693_4 ( .OUT(na8693_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8693_6 ( .RAM_O2(na8693_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8693_2), .COMP_OUT(1'b0) );
// C_AND////      x60y30     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8694_1 ( .OUT(na8694_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8694_6 ( .RAM_O1(na8694_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8694_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y29     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8695_4 ( .OUT(na8695_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8695_6 ( .RAM_O2(na8695_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8695_2), .COMP_OUT(1'b0) );
// C_AND////      x60y29     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8696_1 ( .OUT(na8696_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8696_6 ( .RAM_O1(na8696_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8696_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y28     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8697_4 ( .OUT(na8697_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8697_6 ( .RAM_O2(na8697_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8697_2), .COMP_OUT(1'b0) );
// C_AND////      x60y28     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8698_1 ( .OUT(na8698_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8698_6 ( .RAM_O1(na8698_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8698_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y27     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8699_4 ( .OUT(na8699_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8699_6 ( .RAM_O2(na8699_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8699_2), .COMP_OUT(1'b0) );
// C_AND////      x60y27     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8700_1 ( .OUT(na8700_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8700_6 ( .RAM_O1(na8700_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8700_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y26     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8701_4 ( .OUT(na8701_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8701_6 ( .RAM_O2(na8701_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8701_2), .COMP_OUT(1'b0) );
// C_AND////      x60y26     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8702_1 ( .OUT(na8702_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8702_6 ( .RAM_O1(na8702_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8702_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y25     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8703_4 ( .OUT(na8703_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8703_6 ( .RAM_O2(na8703_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8703_2), .COMP_OUT(1'b0) );
// C_AND////      x60y25     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8704_1 ( .OUT(na8704_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8704_6 ( .RAM_O1(na8704_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8704_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y20     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8705_1 ( .OUT(na8705_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8705_6 ( .RAM_O1(na8705_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8705_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y19     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8706_1 ( .OUT(na8706_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8706_6 ( .RAM_O1(na8706_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8706_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8707_4 ( .OUT(na8707_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8707_6 ( .RAM_O2(na8707_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8707_2), .COMP_OUT(1'b0) );
// C_AND////      x69y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8708_1 ( .OUT(na8708_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8708_6 ( .RAM_O1(na8708_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8708_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8709_4 ( .OUT(na8709_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8709_6 ( .RAM_O2(na8709_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8709_2), .COMP_OUT(1'b0) );
// C_AND////      x69y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8710_1 ( .OUT(na8710_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8710_6 ( .RAM_O1(na8710_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8710_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y28     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8711_1 ( .OUT(na8711_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8711_6 ( .RAM_O1(na8711_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8711_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x69y27     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8712_1 ( .OUT(na8712_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8712_6 ( .RAM_O1(na8712_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8712_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y26     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8713_4 ( .OUT(na8713_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8713_6 ( .RAM_O2(na8713_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8713_2), .COMP_OUT(1'b0) );
// C_AND////      x69y26     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8714_1 ( .OUT(na8714_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8714_6 ( .RAM_O1(na8714_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8714_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y25     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8715_4 ( .OUT(na8715_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8715_6 ( .RAM_O2(na8715_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8715_2), .COMP_OUT(1'b0) );
// C_AND////      x69y25     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8716_1 ( .OUT(na8716_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8716_6 ( .RAM_O1(na8716_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8716_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y32     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8717_4 ( .OUT(na8717_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8717_5 ( .OUT(na8717_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8717_6 ( .RAM_O2(na8717_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8717_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y32     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8718_1 ( .OUT(na8718_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8718_2 ( .OUT(na8718_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8718_6 ( .RAM_O1(na8718_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8718_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y31     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8719_4 ( .OUT(na8719_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8719_5 ( .OUT(na8719_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8719_6 ( .RAM_O2(na8719_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8719_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y31     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8720_1 ( .OUT(na8720_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8720_2 ( .OUT(na8720_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8720_6 ( .RAM_O1(na8720_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8720_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y32     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8721_4 ( .OUT(na8721_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8721_5 ( .OUT(na8721_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8721_6 ( .RAM_O2(na8721_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8721_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y32     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8722_1 ( .OUT(na8722_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8722_2 ( .OUT(na8722_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8722_6 ( .RAM_O1(na8722_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8722_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y31     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8723_4 ( .OUT(na8723_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8723_5 ( .OUT(na8723_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8723_6 ( .RAM_O2(na8723_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8723_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y31     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8724_1 ( .OUT(na8724_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8724_2 ( .OUT(na8724_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8724_6 ( .RAM_O1(na8724_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8724_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y30     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8725_4 ( .OUT(na8725_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8725_5 ( .OUT(na8725_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8725_6 ( .RAM_O2(na8725_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8725_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y30     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8726_1 ( .OUT(na8726_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8726_2 ( .OUT(na8726_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8726_6 ( .RAM_O1(na8726_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8726_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y29     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8727_4 ( .OUT(na8727_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8727_5 ( .OUT(na8727_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8727_6 ( .RAM_O2(na8727_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8727_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y29     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8728_1 ( .OUT(na8728_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8728_2 ( .OUT(na8728_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8728_6 ( .RAM_O1(na8728_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8728_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y28     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8729_4 ( .OUT(na8729_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8729_5 ( .OUT(na8729_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8729_6 ( .RAM_O2(na8729_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8729_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y28     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8730_1 ( .OUT(na8730_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8730_2 ( .OUT(na8730_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8730_6 ( .RAM_O1(na8730_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8730_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y27     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8731_4 ( .OUT(na8731_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8731_5 ( .OUT(na8731_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8731_6 ( .RAM_O2(na8731_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8731_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y27     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8732_1 ( .OUT(na8732_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8732_2 ( .OUT(na8732_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8732_6 ( .RAM_O1(na8732_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8732_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y26     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8733_4 ( .OUT(na8733_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8733_5 ( .OUT(na8733_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8733_6 ( .RAM_O2(na8733_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8733_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y26     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8734_1 ( .OUT(na8734_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8734_2 ( .OUT(na8734_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8734_6 ( .RAM_O1(na8734_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8734_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y25     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8735_4 ( .OUT(na8735_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8735_5 ( .OUT(na8735_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8735_6 ( .RAM_O2(na8735_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8735_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y25     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8736_1 ( .OUT(na8736_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8736_2 ( .OUT(na8736_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8736_6 ( .RAM_O1(na8736_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8736_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y24     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8737_4 ( .OUT(na8737_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8737_5 ( .OUT(na8737_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8737_6 ( .RAM_O2(na8737_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8737_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y24     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8738_1 ( .OUT(na8738_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8738_2 ( .OUT(na8738_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8738_6 ( .RAM_O1(na8738_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8738_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y23     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8739_4 ( .OUT(na8739_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8739_5 ( .OUT(na8739_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8739_6 ( .RAM_O2(na8739_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8739_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y23     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8740_1 ( .OUT(na8740_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8740_2 ( .OUT(na8740_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8740_6 ( .RAM_O1(na8740_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8740_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y24     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8741_4 ( .OUT(na8741_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8741_5 ( .OUT(na8741_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8741_6 ( .RAM_O2(na8741_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8741_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y24     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8742_1 ( .OUT(na8742_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8742_2 ( .OUT(na8742_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8742_6 ( .RAM_O1(na8742_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8742_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y23     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8743_4 ( .OUT(na8743_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8743_5 ( .OUT(na8743_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8743_6 ( .RAM_O2(na8743_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8743_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y23     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8744_1 ( .OUT(na8744_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8744_2 ( .OUT(na8744_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8744_6 ( .RAM_O1(na8744_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8744_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y22     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8745_4 ( .OUT(na8745_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8745_5 ( .OUT(na8745_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8745_6 ( .RAM_O2(na8745_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8745_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y22     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8746_1 ( .OUT(na8746_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8746_2 ( .OUT(na8746_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8746_6 ( .RAM_O1(na8746_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8746_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y21     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8747_4 ( .OUT(na8747_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8747_5 ( .OUT(na8747_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8747_6 ( .RAM_O2(na8747_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8747_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y21     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8748_1 ( .OUT(na8748_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8748_2 ( .OUT(na8748_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8748_6 ( .RAM_O1(na8748_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8748_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y20     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8749_4 ( .OUT(na8749_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8749_5 ( .OUT(na8749_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8749_6 ( .RAM_O2(na8749_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8749_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y20     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8750_1 ( .OUT(na8750_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8750_2 ( .OUT(na8750_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8750_6 ( .RAM_O1(na8750_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8750_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y19     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8751_4 ( .OUT(na8751_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8751_5 ( .OUT(na8751_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8751_6 ( .RAM_O2(na8751_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8751_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y19     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8752_1 ( .OUT(na8752_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8752_2 ( .OUT(na8752_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8752_6 ( .RAM_O1(na8752_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8752_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y18     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8753_4 ( .OUT(na8753_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8753_5 ( .OUT(na8753_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8753_6 ( .RAM_O2(na8753_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8753_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y18     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8754_1 ( .OUT(na8754_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8754_2 ( .OUT(na8754_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8754_6 ( .RAM_O1(na8754_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8754_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y17     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8755_4 ( .OUT(na8755_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8755_5 ( .OUT(na8755_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8755_6 ( .RAM_O2(na8755_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8755_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y17     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8756_1 ( .OUT(na8756_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8756_2 ( .OUT(na8756_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6653_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8756_6 ( .RAM_O1(na8756_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8756_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y32     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8757_4 ( .OUT(na8757_2), .IN1(1'b1), .IN2(na2891_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8757_6 ( .RAM_O2(na8757_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8757_2), .COMP_OUT(1'b0) );
// C_AND////      x61y32     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8758_1 ( .OUT(na8758_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2891_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8758_6 ( .RAM_O1(na8758_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8758_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y31     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8759_4 ( .OUT(na8759_2), .IN1(1'b1), .IN2(na2891_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8759_6 ( .RAM_O2(na8759_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8759_2), .COMP_OUT(1'b0) );
// C_AND////      x61y31     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8760_1 ( .OUT(na8760_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2891_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8760_6 ( .RAM_O1(na8760_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8760_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y32     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8761_4 ( .OUT(na8761_2), .IN1(1'b1), .IN2(na2891_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8761_6 ( .RAM_O2(na8761_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8761_2), .COMP_OUT(1'b0) );
// C_AND////      x63y32     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8762_1 ( .OUT(na8762_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2891_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8762_6 ( .RAM_O1(na8762_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8762_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y31     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8763_4 ( .OUT(na8763_2), .IN1(1'b1), .IN2(na2891_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8763_6 ( .RAM_O2(na8763_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8763_2), .COMP_OUT(1'b0) );
// C_AND////      x63y31     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8764_1 ( .OUT(na8764_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2891_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8764_6 ( .RAM_O1(na8764_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8764_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y30     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8765_4 ( .OUT(na8765_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8765_6 ( .RAM_O2(na8765_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8765_2), .COMP_OUT(1'b0) );
// C_AND////      x63y30     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8766_1 ( .OUT(na8766_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8766_6 ( .RAM_O1(na8766_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8766_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y29     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8767_4 ( .OUT(na8767_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8767_6 ( .RAM_O2(na8767_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8767_2), .COMP_OUT(1'b0) );
// C_AND////      x63y29     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8768_1 ( .OUT(na8768_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8768_6 ( .RAM_O1(na8768_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8768_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y28     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8769_4 ( .OUT(na8769_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8769_6 ( .RAM_O2(na8769_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8769_2), .COMP_OUT(1'b0) );
// C_AND////      x63y28     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8770_1 ( .OUT(na8770_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8770_6 ( .RAM_O1(na8770_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8770_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y27     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8771_4 ( .OUT(na8771_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2890_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8771_6 ( .RAM_O2(na8771_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8771_2), .COMP_OUT(1'b0) );
// C_AND////      x63y27     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8772_1 ( .OUT(na8772_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2890_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8772_6 ( .RAM_O1(na8772_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8772_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y26     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8773_4 ( .OUT(na8773_2), .IN1(na2888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8773_6 ( .RAM_O2(na8773_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8773_2), .COMP_OUT(1'b0) );
// C_AND////      x63y26     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8774_1 ( .OUT(na8774_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2888_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8774_6 ( .RAM_O1(na8774_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8774_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y25     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8775_4 ( .OUT(na8775_2), .IN1(na2888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8775_6 ( .RAM_O2(na8775_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8775_2), .COMP_OUT(1'b0) );
// C_AND////      x63y25     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8776_1 ( .OUT(na8776_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2888_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8776_6 ( .RAM_O1(na8776_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8776_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y24     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8777_4 ( .OUT(na8777_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2863_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8777_6 ( .RAM_O2(na8777_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8777_2), .COMP_OUT(1'b0) );
// C_AND////      x61y24     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8778_1 ( .OUT(na8778_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2863_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8778_6 ( .RAM_O1(na8778_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8778_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y23     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8779_4 ( .OUT(na8779_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2863_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8779_6 ( .RAM_O2(na8779_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8779_2), .COMP_OUT(1'b0) );
// C_AND////      x61y23     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8780_1 ( .OUT(na8780_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2863_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8780_6 ( .RAM_O1(na8780_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8780_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y24     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8781_4 ( .OUT(na8781_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2862_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8781_6 ( .RAM_O2(na8781_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8781_2), .COMP_OUT(1'b0) );
// C_AND////      x63y24     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8782_1 ( .OUT(na8782_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2862_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8782_6 ( .RAM_O1(na8782_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8782_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y23     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8783_4 ( .OUT(na8783_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2862_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8783_6 ( .RAM_O2(na8783_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8783_2), .COMP_OUT(1'b0) );
// C_AND////      x63y23     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8784_1 ( .OUT(na8784_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2862_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8784_6 ( .RAM_O1(na8784_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8784_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y22     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8785_4 ( .OUT(na8785_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2862_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8785_6 ( .RAM_O2(na8785_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8785_2), .COMP_OUT(1'b0) );
// C_AND////      x63y22     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8786_1 ( .OUT(na8786_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2862_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8786_6 ( .RAM_O1(na8786_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8786_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y21     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8787_4 ( .OUT(na8787_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2862_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8787_6 ( .RAM_O2(na8787_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8787_2), .COMP_OUT(1'b0) );
// C_AND////      x63y21     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8788_1 ( .OUT(na8788_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2862_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8788_6 ( .RAM_O1(na8788_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8788_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y20     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8789_4 ( .OUT(na8789_2), .IN1(1'b1), .IN2(na2861_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8789_6 ( .RAM_O2(na8789_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8789_2), .COMP_OUT(1'b0) );
// C_AND////      x63y20     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8790_1 ( .OUT(na8790_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2861_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8790_6 ( .RAM_O1(na8790_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8790_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y19     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8791_4 ( .OUT(na8791_2), .IN1(1'b1), .IN2(na2861_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8791_6 ( .RAM_O2(na8791_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8791_2), .COMP_OUT(1'b0) );
// C_AND////      x63y19     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8792_1 ( .OUT(na8792_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2861_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8792_6 ( .RAM_O1(na8792_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8792_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y18     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8793_4 ( .OUT(na8793_2), .IN1(1'b1), .IN2(na2861_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8793_6 ( .RAM_O2(na8793_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8793_2), .COMP_OUT(1'b0) );
// C_AND////      x63y18     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8794_1 ( .OUT(na8794_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2861_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8794_6 ( .RAM_O1(na8794_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8794_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y17     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8795_4 ( .OUT(na8795_2), .IN1(1'b1), .IN2(na2861_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8795_6 ( .RAM_O2(na8795_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8795_2), .COMP_OUT(1'b0) );
// C_AND////      x63y17     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8796_1 ( .OUT(na8796_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2861_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8796_6 ( .RAM_O1(na8796_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8796_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x35y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8797_1 ( .OUT(na8797_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8797_6 ( .RAM_O1(na8797_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8797_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y81     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8798_4 ( .OUT(na8798_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3215_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8798_6 ( .RAM_O2(na8798_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8798_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y88     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8799_4 ( .OUT(na8799_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8799_6 ( .RAM_O2(na8799_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8799_2), .COMP_OUT(1'b0) );
// C_AND////      x28y88     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8800_1 ( .OUT(na8800_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8800_6 ( .RAM_O1(na8800_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8800_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y87     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8801_4 ( .OUT(na8801_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8801_6 ( .RAM_O2(na8801_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8801_2), .COMP_OUT(1'b0) );
// C_AND////      x28y87     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8802_1 ( .OUT(na8802_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8802_6 ( .RAM_O1(na8802_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8802_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y86     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8803_4 ( .OUT(na8803_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8803_6 ( .RAM_O2(na8803_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8803_2), .COMP_OUT(1'b0) );
// C_AND////      x28y86     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8804_1 ( .OUT(na8804_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8804_6 ( .RAM_O1(na8804_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8804_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y85     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8805_4 ( .OUT(na8805_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8805_6 ( .RAM_O2(na8805_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8805_2), .COMP_OUT(1'b0) );
// C_AND////      x28y85     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8806_1 ( .OUT(na8806_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8806_6 ( .RAM_O1(na8806_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8806_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y84     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8807_4 ( .OUT(na8807_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8807_6 ( .RAM_O2(na8807_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8807_2), .COMP_OUT(1'b0) );
// C_AND////      x28y84     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8808_1 ( .OUT(na8808_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8808_6 ( .RAM_O1(na8808_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8808_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y83     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8809_4 ( .OUT(na8809_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8809_6 ( .RAM_O2(na8809_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8809_2), .COMP_OUT(1'b0) );
// C_AND////      x28y83     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8810_1 ( .OUT(na8810_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8810_6 ( .RAM_O1(na8810_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8810_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y82     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8811_4 ( .OUT(na8811_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8811_6 ( .RAM_O2(na8811_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8811_2), .COMP_OUT(1'b0) );
// C_AND////      x28y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8812_1 ( .OUT(na8812_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8812_6 ( .RAM_O1(na8812_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8812_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8813_4 ( .OUT(na8813_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8813_6 ( .RAM_O2(na8813_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8813_2), .COMP_OUT(1'b0) );
// C_AND////      x28y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8814_1 ( .OUT(na8814_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8814_6 ( .RAM_O1(na8814_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8814_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x37y84     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8815_1 ( .OUT(na8815_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8815_6 ( .RAM_O1(na8815_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8815_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x37y83     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8816_1 ( .OUT(na8816_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8816_6 ( .RAM_O1(na8816_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8816_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y82     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8817_4 ( .OUT(na8817_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8817_6 ( .RAM_O2(na8817_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8817_2), .COMP_OUT(1'b0) );
// C_AND////      x37y82     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8818_1 ( .OUT(na8818_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8818_6 ( .RAM_O1(na8818_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8818_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y81     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8819_4 ( .OUT(na8819_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8819_6 ( .RAM_O2(na8819_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8819_2), .COMP_OUT(1'b0) );
// C_AND////      x37y81     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8820_1 ( .OUT(na8820_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8820_6 ( .RAM_O1(na8820_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8820_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x30y88     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8821_4 ( .OUT(na8821_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8821_5 ( .OUT(na8821_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8821_6 ( .RAM_O2(na8821_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8821_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x30y88     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8822_1 ( .OUT(na8822_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8822_2 ( .OUT(na8822_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8822_6 ( .RAM_O1(na8822_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8822_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x30y87     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8823_4 ( .OUT(na8823_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8823_5 ( .OUT(na8823_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8823_6 ( .RAM_O2(na8823_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8823_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x30y87     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8824_1 ( .OUT(na8824_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8824_2 ( .OUT(na8824_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8824_6 ( .RAM_O1(na8824_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8824_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y88     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8825_4 ( .OUT(na8825_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8825_5 ( .OUT(na8825_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8825_6 ( .RAM_O2(na8825_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8825_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y88     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8826_1 ( .OUT(na8826_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8826_2 ( .OUT(na8826_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8826_6 ( .RAM_O1(na8826_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8826_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y87     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8827_4 ( .OUT(na8827_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8827_5 ( .OUT(na8827_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8827_6 ( .RAM_O2(na8827_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8827_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y87     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8828_1 ( .OUT(na8828_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8828_2 ( .OUT(na8828_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8828_6 ( .RAM_O1(na8828_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8828_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y86     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8829_4 ( .OUT(na8829_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8829_5 ( .OUT(na8829_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8829_6 ( .RAM_O2(na8829_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8829_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y86     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8830_1 ( .OUT(na8830_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8830_2 ( .OUT(na8830_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8830_6 ( .RAM_O1(na8830_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8830_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y85     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8831_4 ( .OUT(na8831_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8831_5 ( .OUT(na8831_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8831_6 ( .RAM_O2(na8831_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8831_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y85     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8832_1 ( .OUT(na8832_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8832_2 ( .OUT(na8832_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8832_6 ( .RAM_O1(na8832_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8832_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y84     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8833_4 ( .OUT(na8833_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8833_5 ( .OUT(na8833_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8833_6 ( .RAM_O2(na8833_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8833_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y84     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8834_1 ( .OUT(na8834_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8834_2 ( .OUT(na8834_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8834_6 ( .RAM_O1(na8834_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8834_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y83     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8835_4 ( .OUT(na8835_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8835_5 ( .OUT(na8835_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8835_6 ( .RAM_O2(na8835_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8835_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y83     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8836_1 ( .OUT(na8836_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8836_2 ( .OUT(na8836_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8836_6 ( .RAM_O1(na8836_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8836_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y82     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8837_4 ( .OUT(na8837_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8837_5 ( .OUT(na8837_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8837_6 ( .RAM_O2(na8837_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8837_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y82     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8838_1 ( .OUT(na8838_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8838_2 ( .OUT(na8838_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8838_6 ( .RAM_O1(na8838_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8838_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x32y81     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8839_4 ( .OUT(na8839_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8839_5 ( .OUT(na8839_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8839_6 ( .RAM_O2(na8839_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8839_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x32y81     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8840_1 ( .OUT(na8840_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8840_2 ( .OUT(na8840_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6655_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8840_6 ( .RAM_O1(na8840_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8840_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y88     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8841_4 ( .OUT(na8841_2), .IN1(1'b1), .IN2(na2870_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8841_6 ( .RAM_O2(na8841_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8841_2), .COMP_OUT(1'b0) );
// C_AND////      x29y88     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8842_1 ( .OUT(na8842_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2870_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8842_6 ( .RAM_O1(na8842_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8842_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y87     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8843_4 ( .OUT(na8843_2), .IN1(1'b1), .IN2(na2870_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8843_6 ( .RAM_O2(na8843_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8843_2), .COMP_OUT(1'b0) );
// C_AND////      x29y87     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8844_1 ( .OUT(na8844_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2870_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8844_6 ( .RAM_O1(na8844_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8844_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y88     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8845_4 ( .OUT(na8845_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2868_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8845_6 ( .RAM_O2(na8845_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8845_2), .COMP_OUT(1'b0) );
// C_AND////      x31y88     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8846_1 ( .OUT(na8846_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2868_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8846_6 ( .RAM_O1(na8846_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8846_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y87     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8847_4 ( .OUT(na8847_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2868_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8847_6 ( .RAM_O2(na8847_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8847_2), .COMP_OUT(1'b0) );
// C_AND////      x31y87     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8848_1 ( .OUT(na8848_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2868_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8848_6 ( .RAM_O1(na8848_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8848_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y86     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8849_4 ( .OUT(na8849_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2868_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8849_6 ( .RAM_O2(na8849_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8849_2), .COMP_OUT(1'b0) );
// C_AND////      x31y86     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8850_1 ( .OUT(na8850_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2868_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8850_6 ( .RAM_O1(na8850_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8850_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y85     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8851_4 ( .OUT(na8851_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2868_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8851_6 ( .RAM_O2(na8851_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8851_2), .COMP_OUT(1'b0) );
// C_AND////      x31y85     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8852_1 ( .OUT(na8852_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2868_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8852_6 ( .RAM_O1(na8852_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8852_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y84     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8853_4 ( .OUT(na8853_2), .IN1(na2867_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8853_6 ( .RAM_O2(na8853_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8853_2), .COMP_OUT(1'b0) );
// C_AND////      x31y84     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8854_1 ( .OUT(na8854_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2867_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8854_6 ( .RAM_O1(na8854_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8854_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y83     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8855_4 ( .OUT(na8855_2), .IN1(na2867_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8855_6 ( .RAM_O2(na8855_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8855_2), .COMP_OUT(1'b0) );
// C_AND////      x31y83     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8856_1 ( .OUT(na8856_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2867_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8856_6 ( .RAM_O1(na8856_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8856_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y82     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8857_4 ( .OUT(na8857_2), .IN1(na2867_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8857_6 ( .RAM_O2(na8857_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8857_2), .COMP_OUT(1'b0) );
// C_AND////      x31y82     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8858_1 ( .OUT(na8858_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2867_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8858_6 ( .RAM_O1(na8858_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8858_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y81     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8859_4 ( .OUT(na8859_2), .IN1(na2867_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8859_6 ( .RAM_O2(na8859_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8859_2), .COMP_OUT(1'b0) );
// C_AND////      x31y81     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8860_1 ( .OUT(na8860_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2867_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8860_6 ( .RAM_O1(na8860_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8860_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x99y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8861_1 ( .OUT(na8861_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8861_6 ( .RAM_O1(na8861_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8861_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x99y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8862_1 ( .OUT(na8862_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8862_6 ( .RAM_O1(na8862_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8862_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x91y57     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8863_4 ( .OUT(na8863_2), .IN1(1'b1), .IN2(na3289_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8863_6 ( .RAM_O2(na8863_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8863_2), .COMP_OUT(1'b0) );
// C_///AND/      x91y49     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8864_4 ( .OUT(na8864_2), .IN1(1'b1), .IN2(na3304_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8864_6 ( .RAM_O2(na8864_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8864_2), .COMP_OUT(1'b0) );
// C_///AND/      x92y56     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8865_4 ( .OUT(na8865_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8865_6 ( .RAM_O2(na8865_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8865_2), .COMP_OUT(1'b0) );
// C_AND////      x92y56     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8866_1 ( .OUT(na8866_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8866_6 ( .RAM_O1(na8866_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8866_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y55     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8867_4 ( .OUT(na8867_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8867_6 ( .RAM_O2(na8867_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8867_2), .COMP_OUT(1'b0) );
// C_AND////      x92y55     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8868_1 ( .OUT(na8868_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8868_6 ( .RAM_O1(na8868_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8868_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y54     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8869_4 ( .OUT(na8869_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8869_6 ( .RAM_O2(na8869_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8869_2), .COMP_OUT(1'b0) );
// C_AND////      x92y54     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8870_1 ( .OUT(na8870_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8870_6 ( .RAM_O1(na8870_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8870_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y53     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8871_4 ( .OUT(na8871_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8871_6 ( .RAM_O2(na8871_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8871_2), .COMP_OUT(1'b0) );
// C_AND////      x92y53     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8872_1 ( .OUT(na8872_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8872_6 ( .RAM_O1(na8872_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8872_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y52     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8873_4 ( .OUT(na8873_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8873_6 ( .RAM_O2(na8873_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8873_2), .COMP_OUT(1'b0) );
// C_AND////      x92y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8874_1 ( .OUT(na8874_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8874_6 ( .RAM_O1(na8874_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8874_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y51     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8875_4 ( .OUT(na8875_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8875_6 ( .RAM_O2(na8875_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8875_2), .COMP_OUT(1'b0) );
// C_AND////      x92y51     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8876_1 ( .OUT(na8876_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8876_6 ( .RAM_O1(na8876_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8876_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8877_4 ( .OUT(na8877_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8877_6 ( .RAM_O2(na8877_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8877_2), .COMP_OUT(1'b0) );
// C_AND////      x92y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8878_1 ( .OUT(na8878_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8878_6 ( .RAM_O1(na8878_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8878_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8879_4 ( .OUT(na8879_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8879_6 ( .RAM_O2(na8879_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8879_2), .COMP_OUT(1'b0) );
// C_AND////      x92y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8880_1 ( .OUT(na8880_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8880_6 ( .RAM_O1(na8880_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8880_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y64     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8881_4 ( .OUT(na8881_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8881_6 ( .RAM_O2(na8881_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8881_2), .COMP_OUT(1'b0) );
// C_AND////      x92y64     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8882_1 ( .OUT(na8882_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na86_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8882_6 ( .RAM_O1(na8882_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8882_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y63     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8883_4 ( .OUT(na8883_2), .IN1(1'b1), .IN2(na85_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8883_6 ( .RAM_O2(na8883_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8883_2), .COMP_OUT(1'b0) );
// C_AND////      x92y63     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8884_1 ( .OUT(na8884_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na84_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8884_6 ( .RAM_O1(na8884_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8884_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y62     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8885_4 ( .OUT(na8885_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8885_6 ( .RAM_O2(na8885_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8885_2), .COMP_OUT(1'b0) );
// C_AND////      x92y62     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8886_1 ( .OUT(na8886_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na35_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8886_6 ( .RAM_O1(na8886_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8886_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y61     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8887_4 ( .OUT(na8887_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na37_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8887_6 ( .RAM_O2(na8887_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8887_2), .COMP_OUT(1'b0) );
// C_AND////      x92y61     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8888_1 ( .OUT(na8888_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8888_6 ( .RAM_O1(na8888_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8888_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y60     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8889_4 ( .OUT(na8889_2), .IN1(1'b1), .IN2(1'b1), .IN3(na66_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8889_6 ( .RAM_O2(na8889_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8889_2), .COMP_OUT(1'b0) );
// C_AND////      x92y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8890_1 ( .OUT(na8890_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8890_6 ( .RAM_O1(na8890_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8890_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y59     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8891_4 ( .OUT(na8891_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8891_6 ( .RAM_O2(na8891_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8891_2), .COMP_OUT(1'b0) );
// C_AND////      x92y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8892_1 ( .OUT(na8892_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8892_6 ( .RAM_O1(na8892_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8892_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8893_4 ( .OUT(na8893_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8893_6 ( .RAM_O2(na8893_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8893_2), .COMP_OUT(1'b0) );
// C_AND////      x92y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8894_1 ( .OUT(na8894_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8894_6 ( .RAM_O1(na8894_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8894_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x92y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8895_4 ( .OUT(na8895_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8895_6 ( .RAM_O2(na8895_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8895_2), .COMP_OUT(1'b0) );
// C_AND////      x92y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8896_1 ( .OUT(na8896_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8896_6 ( .RAM_O1(na8896_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8896_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x101y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8897_1 ( .OUT(na8897_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8897_6 ( .RAM_O1(na8897_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8897_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x101y51     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8898_1 ( .OUT(na8898_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8898_6 ( .RAM_O1(na8898_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8898_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8899_4 ( .OUT(na8899_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8899_6 ( .RAM_O2(na8899_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8899_2), .COMP_OUT(1'b0) );
// C_AND////      x101y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8900_1 ( .OUT(na8900_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8900_6 ( .RAM_O1(na8900_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8900_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8901_4 ( .OUT(na8901_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8901_6 ( .RAM_O2(na8901_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8901_2), .COMP_OUT(1'b0) );
// C_AND////      x101y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8902_1 ( .OUT(na8902_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8902_6 ( .RAM_O1(na8902_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8902_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x101y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8903_1 ( .OUT(na8903_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8903_6 ( .RAM_O1(na8903_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8903_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x101y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8904_1 ( .OUT(na8904_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8904_6 ( .RAM_O1(na8904_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8904_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8905_4 ( .OUT(na8905_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8905_6 ( .RAM_O2(na8905_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8905_2), .COMP_OUT(1'b0) );
// C_AND////      x101y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8906_1 ( .OUT(na8906_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8906_6 ( .RAM_O1(na8906_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8906_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x101y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8907_4 ( .OUT(na8907_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8907_6 ( .RAM_O2(na8907_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8907_2), .COMP_OUT(1'b0) );
// C_AND////      x101y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8908_1 ( .OUT(na8908_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8908_6 ( .RAM_O1(na8908_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8908_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x94y64     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8909_4 ( .OUT(na8909_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2551_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8909_5 ( .OUT(na8909_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8909_6 ( .RAM_O2(na8909_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8909_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x94y64     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8910_1 ( .OUT(na8910_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2550_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8910_2 ( .OUT(na8910_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8910_6 ( .RAM_O1(na8910_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8910_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x94y63     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8911_4 ( .OUT(na8911_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8911_5 ( .OUT(na8911_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8911_6 ( .RAM_O2(na8911_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8911_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x94y63     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8912_1 ( .OUT(na8912_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8912_2 ( .OUT(na8912_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8912_6 ( .RAM_O1(na8912_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8912_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y64     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8913_4 ( .OUT(na8913_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2547_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8913_5 ( .OUT(na8913_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8913_6 ( .RAM_O2(na8913_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8913_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y64     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8914_1 ( .OUT(na8914_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2546_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8914_2 ( .OUT(na8914_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8914_6 ( .RAM_O1(na8914_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8914_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y63     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8915_4 ( .OUT(na8915_2_i), .IN1(1'b1), .IN2(na2545_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8915_5 ( .OUT(na8915_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8915_6 ( .RAM_O2(na8915_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8915_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y63     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8916_1 ( .OUT(na8916_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2544_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8916_2 ( .OUT(na8916_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8916_6 ( .RAM_O1(na8916_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8916_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y62     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8917_4 ( .OUT(na8917_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8917_5 ( .OUT(na8917_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8917_6 ( .RAM_O2(na8917_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8917_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y62     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8918_1 ( .OUT(na8918_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2542_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8918_2 ( .OUT(na8918_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8918_6 ( .RAM_O1(na8918_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8918_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y61     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8919_4 ( .OUT(na8919_2_i), .IN1(na2541_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8919_5 ( .OUT(na8919_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8919_6 ( .RAM_O2(na8919_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8919_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y61     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8920_1 ( .OUT(na8920_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2540_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8920_2 ( .OUT(na8920_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8920_6 ( .RAM_O1(na8920_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8920_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y60     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8921_4 ( .OUT(na8921_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8921_5 ( .OUT(na8921_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8921_6 ( .RAM_O2(na8921_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8921_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y60     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8922_1 ( .OUT(na8922_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8922_2 ( .OUT(na8922_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8922_6 ( .RAM_O1(na8922_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8922_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y59     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8923_4 ( .OUT(na8923_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8923_5 ( .OUT(na8923_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8923_6 ( .RAM_O2(na8923_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8923_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y59     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8924_1 ( .OUT(na8924_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8924_2 ( .OUT(na8924_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8924_6 ( .RAM_O1(na8924_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8924_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y58     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8925_4 ( .OUT(na8925_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8925_5 ( .OUT(na8925_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8925_6 ( .RAM_O2(na8925_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8925_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y58     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8926_1 ( .OUT(na8926_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8926_2 ( .OUT(na8926_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8926_6 ( .RAM_O1(na8926_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8926_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y57     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8927_4 ( .OUT(na8927_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8927_5 ( .OUT(na8927_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8927_6 ( .RAM_O2(na8927_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8927_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y57     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8928_1 ( .OUT(na8928_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8928_2 ( .OUT(na8928_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8928_6 ( .RAM_O1(na8928_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8928_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x94y56     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8929_4 ( .OUT(na8929_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8929_5 ( .OUT(na8929_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8929_6 ( .RAM_O2(na8929_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8929_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x94y56     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8930_1 ( .OUT(na8930_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2538_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8930_2 ( .OUT(na8930_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8930_6 ( .RAM_O1(na8930_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8930_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x94y55     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8931_4 ( .OUT(na8931_2_i), .IN1(na2537_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8931_5 ( .OUT(na8931_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8931_6 ( .RAM_O2(na8931_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8931_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x94y55     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8932_1 ( .OUT(na8932_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2536_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8932_2 ( .OUT(na8932_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8932_6 ( .RAM_O1(na8932_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8932_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y56     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8933_4 ( .OUT(na8933_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8933_5 ( .OUT(na8933_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8933_6 ( .RAM_O2(na8933_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8933_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y56     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8934_1 ( .OUT(na8934_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8934_2 ( .OUT(na8934_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8934_6 ( .RAM_O1(na8934_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8934_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y55     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8935_4 ( .OUT(na8935_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8935_5 ( .OUT(na8935_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8935_6 ( .RAM_O2(na8935_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8935_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y55     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8936_1 ( .OUT(na8936_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2528_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8936_2 ( .OUT(na8936_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8936_6 ( .RAM_O1(na8936_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8936_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y54     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8937_4 ( .OUT(na8937_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2526_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8937_5 ( .OUT(na8937_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8937_6 ( .RAM_O2(na8937_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8937_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y54     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8938_1 ( .OUT(na8938_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2524_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8938_2 ( .OUT(na8938_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8938_6 ( .RAM_O1(na8938_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8938_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y53     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8939_4 ( .OUT(na8939_2_i), .IN1(na2522_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8939_5 ( .OUT(na8939_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8939_6 ( .RAM_O2(na8939_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8939_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y53     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8940_1 ( .OUT(na8940_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2520_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8940_2 ( .OUT(na8940_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8940_6 ( .RAM_O1(na8940_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8940_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y52     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8941_4 ( .OUT(na8941_2_i), .IN1(1'b1), .IN2(na5593_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8941_5 ( .OUT(na8941_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8941_6 ( .RAM_O2(na8941_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8941_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y52     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8942_1 ( .OUT(na8942_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5592_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8942_2 ( .OUT(na8942_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8942_6 ( .RAM_O1(na8942_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8942_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y51     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8943_4 ( .OUT(na8943_2_i), .IN1(na5591_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8943_5 ( .OUT(na8943_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8943_6 ( .RAM_O2(na8943_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8943_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y51     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8944_1 ( .OUT(na8944_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5590_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8944_2 ( .OUT(na8944_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8944_6 ( .RAM_O1(na8944_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8944_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y50     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8945_4 ( .OUT(na8945_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na5589_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8945_5 ( .OUT(na8945_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8945_6 ( .RAM_O2(na8945_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8945_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y50     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8946_1 ( .OUT(na8946_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5588_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8946_2 ( .OUT(na8946_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8946_6 ( .RAM_O1(na8946_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8946_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x96y49     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8947_4 ( .OUT(na8947_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na5587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8947_5 ( .OUT(na8947_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8947_6 ( .RAM_O2(na8947_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8947_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x96y49     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8948_1 ( .OUT(na8948_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na5586_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a8948_2 ( .OUT(na8948_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6657_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8948_6 ( .RAM_O1(na8948_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8948_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y64     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8949_4 ( .OUT(na8949_2), .IN1(na2872_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8949_6 ( .RAM_O2(na8949_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8949_2), .COMP_OUT(1'b0) );
// C_AND////      x93y64     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8950_1 ( .OUT(na8950_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2872_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8950_6 ( .RAM_O1(na8950_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8950_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y63     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8951_4 ( .OUT(na8951_2), .IN1(na2872_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8951_6 ( .RAM_O2(na8951_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8951_2), .COMP_OUT(1'b0) );
// C_AND////      x93y63     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8952_1 ( .OUT(na8952_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2872_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8952_6 ( .RAM_O1(na8952_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8952_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y64     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8953_4 ( .OUT(na8953_2), .IN1(na2872_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8953_6 ( .RAM_O2(na8953_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8953_2), .COMP_OUT(1'b0) );
// C_AND////      x95y64     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8954_1 ( .OUT(na8954_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2872_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8954_6 ( .RAM_O1(na8954_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8954_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y63     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8955_4 ( .OUT(na8955_2), .IN1(na2872_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8955_6 ( .RAM_O2(na8955_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8955_2), .COMP_OUT(1'b0) );
// C_AND////      x95y63     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8956_1 ( .OUT(na8956_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2872_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8956_6 ( .RAM_O1(na8956_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8956_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y62     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8957_4 ( .OUT(na8957_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2871_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8957_6 ( .RAM_O2(na8957_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8957_2), .COMP_OUT(1'b0) );
// C_AND////      x95y62     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8958_1 ( .OUT(na8958_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2871_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8958_6 ( .RAM_O1(na8958_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8958_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y61     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8959_4 ( .OUT(na8959_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2871_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8959_6 ( .RAM_O2(na8959_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8959_2), .COMP_OUT(1'b0) );
// C_AND////      x95y61     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8960_1 ( .OUT(na8960_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2871_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8960_6 ( .RAM_O1(na8960_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8960_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y60     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8961_4 ( .OUT(na8961_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2871_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8961_6 ( .RAM_O2(na8961_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8961_2), .COMP_OUT(1'b0) );
// C_AND////      x95y60     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8962_1 ( .OUT(na8962_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2871_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8962_6 ( .RAM_O1(na8962_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8962_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y59     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8963_4 ( .OUT(na8963_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2871_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8963_6 ( .RAM_O2(na8963_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8963_2), .COMP_OUT(1'b0) );
// C_AND////      x95y59     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8964_1 ( .OUT(na8964_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2871_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8964_6 ( .RAM_O1(na8964_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8964_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y58     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8965_4 ( .OUT(na8965_2), .IN1(1'b1), .IN2(na2870_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8965_6 ( .RAM_O2(na8965_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8965_2), .COMP_OUT(1'b0) );
// C_AND////      x95y58     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8966_1 ( .OUT(na8966_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2870_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8966_6 ( .RAM_O1(na8966_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8966_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y57     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8967_4 ( .OUT(na8967_2), .IN1(1'b1), .IN2(na2870_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8967_6 ( .RAM_O2(na8967_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8967_2), .COMP_OUT(1'b0) );
// C_AND////      x95y57     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8968_1 ( .OUT(na8968_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2870_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8968_6 ( .RAM_O1(na8968_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8968_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y56     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8969_4 ( .OUT(na8969_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2876_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8969_6 ( .RAM_O2(na8969_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8969_2), .COMP_OUT(1'b0) );
// C_AND////      x93y56     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8970_1 ( .OUT(na8970_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2876_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8970_6 ( .RAM_O1(na8970_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8970_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y55     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8971_4 ( .OUT(na8971_2), .IN1(1'b1), .IN2(1'b1), .IN3(na2876_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8971_6 ( .RAM_O2(na8971_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8971_2), .COMP_OUT(1'b0) );
// C_AND////      x93y55     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8972_1 ( .OUT(na8972_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2876_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8972_6 ( .RAM_O1(na8972_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8972_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y56     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8973_4 ( .OUT(na8973_2), .IN1(na2875_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8973_6 ( .RAM_O2(na8973_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8973_2), .COMP_OUT(1'b0) );
// C_AND////      x95y56     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8974_1 ( .OUT(na8974_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2875_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8974_6 ( .RAM_O1(na8974_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8974_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y55     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8975_4 ( .OUT(na8975_2), .IN1(na2875_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8975_6 ( .RAM_O2(na8975_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8975_2), .COMP_OUT(1'b0) );
// C_AND////      x95y55     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8976_1 ( .OUT(na8976_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2875_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8976_6 ( .RAM_O1(na8976_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8976_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y54     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8977_4 ( .OUT(na8977_2), .IN1(na2875_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8977_6 ( .RAM_O2(na8977_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8977_2), .COMP_OUT(1'b0) );
// C_AND////      x95y54     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8978_1 ( .OUT(na8978_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2875_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8978_6 ( .RAM_O1(na8978_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8978_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y53     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8979_4 ( .OUT(na8979_2), .IN1(na2875_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8979_6 ( .RAM_O2(na8979_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8979_2), .COMP_OUT(1'b0) );
// C_AND////      x95y53     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8980_1 ( .OUT(na8980_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2875_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8980_6 ( .RAM_O1(na8980_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8980_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y52     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8981_4 ( .OUT(na8981_2), .IN1(1'b1), .IN2(na2873_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8981_6 ( .RAM_O2(na8981_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8981_2), .COMP_OUT(1'b0) );
// C_AND////      x95y52     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8982_1 ( .OUT(na8982_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2873_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8982_6 ( .RAM_O1(na8982_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8982_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y51     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8983_4 ( .OUT(na8983_2), .IN1(1'b1), .IN2(na2873_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8983_6 ( .RAM_O2(na8983_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8983_2), .COMP_OUT(1'b0) );
// C_AND////      x95y51     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8984_1 ( .OUT(na8984_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2873_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8984_6 ( .RAM_O1(na8984_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8984_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y50     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8985_4 ( .OUT(na8985_2), .IN1(1'b1), .IN2(na2873_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8985_6 ( .RAM_O2(na8985_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8985_2), .COMP_OUT(1'b0) );
// C_AND////      x95y50     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8986_1 ( .OUT(na8986_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2873_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8986_6 ( .RAM_O1(na8986_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8986_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x95y49     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8987_4 ( .OUT(na8987_2), .IN1(1'b1), .IN2(na2873_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8987_6 ( .RAM_O2(na8987_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8987_2), .COMP_OUT(1'b0) );
// C_AND////      x95y49     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8988_1 ( .OUT(na8988_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2873_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8988_6 ( .RAM_O1(na8988_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8988_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x67y58     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8989_1 ( .OUT(na8989_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8989_6 ( .RAM_O1(na8989_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8989_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x67y50     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8990_1 ( .OUT(na8990_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1136_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8990_6 ( .RAM_O1(na8990_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8990_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x59y57     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8991_4 ( .OUT(na8991_2), .IN1(1'b1), .IN2(na1181_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8991_6 ( .RAM_O2(na8991_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8991_2), .COMP_OUT(1'b0) );
// C_///AND/      x59y49     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8992_4 ( .OUT(na8992_2), .IN1(1'b1), .IN2(na1130_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8992_6 ( .RAM_O2(na8992_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8992_2), .COMP_OUT(1'b0) );
// C_///AND/      x60y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8993_4 ( .OUT(na8993_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8993_6 ( .RAM_O2(na8993_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8993_2), .COMP_OUT(1'b0) );
// C_AND////      x60y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8994_1 ( .OUT(na8994_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8994_6 ( .RAM_O1(na8994_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8994_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8995_4 ( .OUT(na8995_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8995_6 ( .RAM_O2(na8995_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8995_2), .COMP_OUT(1'b0) );
// C_AND////      x60y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8996_1 ( .OUT(na8996_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8996_6 ( .RAM_O1(na8996_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8996_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y54     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8997_4 ( .OUT(na8997_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8997_6 ( .RAM_O2(na8997_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8997_2), .COMP_OUT(1'b0) );
// C_AND////      x60y54     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8998_1 ( .OUT(na8998_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8998_6 ( .RAM_O1(na8998_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na8998_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y53     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8999_4 ( .OUT(na8999_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a8999_6 ( .RAM_O2(na8999_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na8999_2), .COMP_OUT(1'b0) );
// C_AND////      x60y53     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9000_1 ( .OUT(na9000_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4135_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9000_6 ( .RAM_O1(na9000_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9000_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y52     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9001_4 ( .OUT(na9001_2), .IN1(1'b1), .IN2(na4134_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9001_6 ( .RAM_O2(na9001_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9001_2), .COMP_OUT(1'b0) );
// C_AND////      x60y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9002_1 ( .OUT(na9002_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9002_6 ( .RAM_O1(na9002_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9002_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y51     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9003_4 ( .OUT(na9003_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4133_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9003_6 ( .RAM_O2(na9003_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9003_2), .COMP_OUT(1'b0) );
// C_AND////      x60y51     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9004_1 ( .OUT(na9004_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4132_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9004_6 ( .RAM_O1(na9004_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9004_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9005_4 ( .OUT(na9005_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9005_6 ( .RAM_O2(na9005_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9005_2), .COMP_OUT(1'b0) );
// C_AND////      x60y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9006_1 ( .OUT(na9006_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9006_6 ( .RAM_O1(na9006_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9006_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9007_4 ( .OUT(na9007_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9007_6 ( .RAM_O2(na9007_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9007_2), .COMP_OUT(1'b0) );
// C_AND////      x60y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9008_1 ( .OUT(na9008_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9008_6 ( .RAM_O1(na9008_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9008_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9009_4 ( .OUT(na9009_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9009_6 ( .RAM_O2(na9009_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9009_2), .COMP_OUT(1'b0) );
// C_AND////      x60y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9010_1 ( .OUT(na9010_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9010_6 ( .RAM_O1(na9010_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9010_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9011_4 ( .OUT(na9011_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9011_6 ( .RAM_O2(na9011_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9011_2), .COMP_OUT(1'b0) );
// C_AND////      x60y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9012_1 ( .OUT(na9012_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9012_6 ( .RAM_O1(na9012_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9012_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9013_4 ( .OUT(na9013_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9013_6 ( .RAM_O2(na9013_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9013_2), .COMP_OUT(1'b0) );
// C_AND////      x60y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9014_1 ( .OUT(na9014_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9014_6 ( .RAM_O1(na9014_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9014_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y61     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9015_4 ( .OUT(na9015_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9015_6 ( .RAM_O2(na9015_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9015_2), .COMP_OUT(1'b0) );
// C_AND////      x60y61     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9016_1 ( .OUT(na9016_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4141_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9016_6 ( .RAM_O1(na9016_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9016_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y60     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9017_4 ( .OUT(na9017_2), .IN1(1'b1), .IN2(1'b1), .IN3(na4140_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9017_6 ( .RAM_O2(na9017_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9017_2), .COMP_OUT(1'b0) );
// C_AND////      x60y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9018_1 ( .OUT(na9018_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9018_6 ( .RAM_O1(na9018_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9018_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y59     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9019_4 ( .OUT(na9019_2), .IN1(na4139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9019_6 ( .RAM_O2(na9019_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9019_2), .COMP_OUT(1'b0) );
// C_AND////      x60y59     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9020_1 ( .OUT(na9020_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4138_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9020_6 ( .RAM_O1(na9020_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9020_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9021_4 ( .OUT(na9021_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9021_6 ( .RAM_O2(na9021_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9021_2), .COMP_OUT(1'b0) );
// C_AND////      x60y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9022_1 ( .OUT(na9022_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9022_6 ( .RAM_O1(na9022_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9022_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9023_4 ( .OUT(na9023_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9023_6 ( .RAM_O2(na9023_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9023_2), .COMP_OUT(1'b0) );
// C_AND////      x60y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9024_1 ( .OUT(na9024_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9024_6 ( .RAM_O1(na9024_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9024_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9025_4 ( .OUT(na9025_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9025_6 ( .RAM_O2(na9025_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9025_2), .COMP_OUT(1'b0) );
// C_AND////      x69y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9026_1 ( .OUT(na9026_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9026_6 ( .RAM_O1(na9026_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9026_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9027_4 ( .OUT(na9027_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9027_6 ( .RAM_O2(na9027_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9027_2), .COMP_OUT(1'b0) );
// C_AND////      x69y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9028_1 ( .OUT(na9028_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9028_6 ( .RAM_O1(na9028_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9028_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y54     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9029_4 ( .OUT(na9029_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9029_6 ( .RAM_O2(na9029_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9029_2), .COMP_OUT(1'b0) );
// C_AND////      x69y54     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9030_1 ( .OUT(na9030_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9030_6 ( .RAM_O1(na9030_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9030_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y53     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9031_4 ( .OUT(na9031_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9031_6 ( .RAM_O2(na9031_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9031_2), .COMP_OUT(1'b0) );
// C_AND////      x69y53     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9032_1 ( .OUT(na9032_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1169_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9032_6 ( .RAM_O1(na9032_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9032_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y52     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9033_4 ( .OUT(na9033_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1170_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9033_6 ( .RAM_O2(na9033_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9033_2), .COMP_OUT(1'b0) );
// C_AND////      x69y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9034_1 ( .OUT(na9034_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9034_6 ( .RAM_O1(na9034_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9034_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y51     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9035_4 ( .OUT(na9035_2), .IN1(na1171_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9035_6 ( .RAM_O2(na9035_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9035_2), .COMP_OUT(1'b0) );
// C_AND////      x69y51     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9036_1 ( .OUT(na9036_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1172_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9036_6 ( .RAM_O1(na9036_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9036_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9037_4 ( .OUT(na9037_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9037_6 ( .RAM_O2(na9037_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9037_2), .COMP_OUT(1'b0) );
// C_AND////      x69y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9038_1 ( .OUT(na9038_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9038_6 ( .RAM_O1(na9038_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9038_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9039_4 ( .OUT(na9039_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9039_6 ( .RAM_O2(na9039_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9039_2), .COMP_OUT(1'b0) );
// C_AND////      x69y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9040_1 ( .OUT(na9040_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9040_6 ( .RAM_O1(na9040_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9040_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9041_4 ( .OUT(na9041_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9041_6 ( .RAM_O2(na9041_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9041_2), .COMP_OUT(1'b0) );
// C_AND////      x69y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9042_1 ( .OUT(na9042_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9042_6 ( .RAM_O1(na9042_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9042_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9043_4 ( .OUT(na9043_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9043_6 ( .RAM_O2(na9043_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9043_2), .COMP_OUT(1'b0) );
// C_AND////      x69y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9044_1 ( .OUT(na9044_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9044_6 ( .RAM_O1(na9044_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9044_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9045_4 ( .OUT(na9045_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9045_6 ( .RAM_O2(na9045_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9045_2), .COMP_OUT(1'b0) );
// C_AND////      x69y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9046_1 ( .OUT(na9046_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9046_6 ( .RAM_O1(na9046_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9046_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y61     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9047_4 ( .OUT(na9047_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9047_6 ( .RAM_O2(na9047_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9047_2), .COMP_OUT(1'b0) );
// C_AND////      x69y61     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9048_1 ( .OUT(na9048_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1219_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9048_6 ( .RAM_O1(na9048_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9048_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y60     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9049_4 ( .OUT(na9049_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1220_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9049_6 ( .RAM_O2(na9049_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9049_2), .COMP_OUT(1'b0) );
// C_AND////      x69y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9050_1 ( .OUT(na9050_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9050_6 ( .RAM_O1(na9050_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9050_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y59     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9051_4 ( .OUT(na9051_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1221_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9051_6 ( .RAM_O2(na9051_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9051_2), .COMP_OUT(1'b0) );
// C_AND////      x69y59     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9052_1 ( .OUT(na9052_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1222_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9052_6 ( .RAM_O1(na9052_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9052_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9053_4 ( .OUT(na9053_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9053_6 ( .RAM_O2(na9053_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9053_2), .COMP_OUT(1'b0) );
// C_AND////      x69y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9054_1 ( .OUT(na9054_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9054_6 ( .RAM_O1(na9054_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9054_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9055_4 ( .OUT(na9055_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9055_6 ( .RAM_O2(na9055_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9055_2), .COMP_OUT(1'b0) );
// C_AND////      x69y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9056_1 ( .OUT(na9056_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9056_6 ( .RAM_O1(na9056_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9056_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x62y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9057_4 ( .OUT(na9057_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9057_6 ( .RAM_O2(na9057_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9057_2), .COMP_OUT(1'b0) );
// C_AND////      x62y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9058_1 ( .OUT(na9058_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9058_6 ( .RAM_O1(na9058_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9058_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x62y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9059_4 ( .OUT(na9059_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9059_6 ( .RAM_O2(na9059_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9059_2), .COMP_OUT(1'b0) );
// C_AND////      x62y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9060_1 ( .OUT(na9060_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9060_6 ( .RAM_O1(na9060_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9060_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9061_4 ( .OUT(na9061_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9061_6 ( .RAM_O2(na9061_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9061_2), .COMP_OUT(1'b0) );
// C_AND////      x64y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9062_1 ( .OUT(na9062_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9062_6 ( .RAM_O1(na9062_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9062_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9063_4 ( .OUT(na9063_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9063_6 ( .RAM_O2(na9063_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9063_2), .COMP_OUT(1'b0) );
// C_AND////      x64y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9064_1 ( .OUT(na9064_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9064_6 ( .RAM_O1(na9064_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9064_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9065_4 ( .OUT(na9065_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9065_6 ( .RAM_O2(na9065_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9065_2), .COMP_OUT(1'b0) );
// C_AND////      x64y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9066_1 ( .OUT(na9066_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9066_6 ( .RAM_O1(na9066_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9066_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y61     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9067_4 ( .OUT(na9067_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9067_6 ( .RAM_O2(na9067_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9067_2), .COMP_OUT(1'b0) );
// C_AND////      x64y61     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9068_1 ( .OUT(na9068_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9068_6 ( .RAM_O1(na9068_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9068_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y60     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9069_4 ( .OUT(na9069_2), .IN1(na419_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9069_6 ( .RAM_O2(na9069_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9069_2), .COMP_OUT(1'b0) );
// C_AND////      x64y60     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9070_1 ( .OUT(na9070_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na418_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9070_6 ( .RAM_O1(na9070_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9070_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y59     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9071_4 ( .OUT(na9071_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na416_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9071_6 ( .RAM_O2(na9071_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9071_2), .COMP_OUT(1'b0) );
// C_AND////      x64y59     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9072_1 ( .OUT(na9072_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na415_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9072_6 ( .RAM_O1(na9072_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9072_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y58     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9073_4 ( .OUT(na9073_2), .IN1(1'b1), .IN2(na414_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9073_6 ( .RAM_O2(na9073_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9073_2), .COMP_OUT(1'b0) );
// C_AND////      x64y58     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9074_1 ( .OUT(na9074_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na413_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9074_6 ( .RAM_O1(na9074_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9074_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y57     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9075_4 ( .OUT(na9075_2), .IN1(na412_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9075_6 ( .RAM_O2(na9075_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9075_2), .COMP_OUT(1'b0) );
// C_AND////      x64y57     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9076_1 ( .OUT(na9076_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na408_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9076_6 ( .RAM_O1(na9076_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9076_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x62y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9077_4 ( .OUT(na9077_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9077_6 ( .RAM_O2(na9077_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9077_2), .COMP_OUT(1'b0) );
// C_AND////      x62y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9078_1 ( .OUT(na9078_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9078_6 ( .RAM_O1(na9078_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9078_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x62y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9079_4 ( .OUT(na9079_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9079_6 ( .RAM_O2(na9079_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9079_2), .COMP_OUT(1'b0) );
// C_AND////      x62y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9080_1 ( .OUT(na9080_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9080_6 ( .RAM_O1(na9080_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9080_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9081_4 ( .OUT(na9081_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9081_6 ( .RAM_O2(na9081_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9081_2), .COMP_OUT(1'b0) );
// C_AND////      x64y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9082_1 ( .OUT(na9082_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9082_6 ( .RAM_O1(na9082_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9082_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9083_4 ( .OUT(na9083_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9083_6 ( .RAM_O2(na9083_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9083_2), .COMP_OUT(1'b0) );
// C_AND////      x64y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9084_1 ( .OUT(na9084_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9084_6 ( .RAM_O1(na9084_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9084_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y54     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9085_4 ( .OUT(na9085_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9085_6 ( .RAM_O2(na9085_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9085_2), .COMP_OUT(1'b0) );
// C_AND////      x64y54     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9086_1 ( .OUT(na9086_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9086_6 ( .RAM_O1(na9086_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9086_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y53     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9087_4 ( .OUT(na9087_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9087_6 ( .RAM_O2(na9087_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9087_2), .COMP_OUT(1'b0) );
// C_AND////      x64y53     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9088_1 ( .OUT(na9088_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9088_6 ( .RAM_O1(na9088_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9088_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y52     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9089_4 ( .OUT(na9089_2), .IN1(1'b1), .IN2(na265_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9089_6 ( .RAM_O2(na9089_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9089_2), .COMP_OUT(1'b0) );
// C_AND////      x64y52     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9090_1 ( .OUT(na9090_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na264_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9090_6 ( .RAM_O1(na9090_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9090_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y51     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9091_4 ( .OUT(na9091_2), .IN1(1'b1), .IN2(1'b1), .IN3(na263_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9091_6 ( .RAM_O2(na9091_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9091_2), .COMP_OUT(1'b0) );
// C_AND////      x64y51     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9092_1 ( .OUT(na9092_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na262_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9092_6 ( .RAM_O1(na9092_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9092_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y50     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9093_4 ( .OUT(na9093_2), .IN1(1'b1), .IN2(1'b1), .IN3(na261_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9093_6 ( .RAM_O2(na9093_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9093_2), .COMP_OUT(1'b0) );
// C_AND////      x64y50     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9094_1 ( .OUT(na9094_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na260_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9094_6 ( .RAM_O1(na9094_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9094_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x64y49     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9095_4 ( .OUT(na9095_2), .IN1(1'b1), .IN2(na259_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9095_6 ( .RAM_O2(na9095_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9095_2), .COMP_OUT(1'b0) );
// C_AND////      x64y49     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9096_1 ( .OUT(na9096_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na159_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9096_6 ( .RAM_O1(na9096_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9096_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9097_4 ( .OUT(na9097_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9097_6 ( .RAM_O2(na9097_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9097_2), .COMP_OUT(1'b0) );
// C_AND////      x61y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9098_1 ( .OUT(na9098_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9098_6 ( .RAM_O1(na9098_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9098_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9099_4 ( .OUT(na9099_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9099_6 ( .RAM_O2(na9099_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9099_2), .COMP_OUT(1'b0) );
// C_AND////      x61y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9100_1 ( .OUT(na9100_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9100_6 ( .RAM_O1(na9100_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9100_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9101_4 ( .OUT(na9101_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9101_6 ( .RAM_O2(na9101_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9101_2), .COMP_OUT(1'b0) );
// C_AND////      x63y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9102_1 ( .OUT(na9102_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9102_6 ( .RAM_O1(na9102_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9102_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9103_4 ( .OUT(na9103_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9103_6 ( .RAM_O2(na9103_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9103_2), .COMP_OUT(1'b0) );
// C_AND////      x63y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9104_1 ( .OUT(na9104_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9104_6 ( .RAM_O1(na9104_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9104_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9105_4 ( .OUT(na9105_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9105_6 ( .RAM_O2(na9105_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9105_2), .COMP_OUT(1'b0) );
// C_AND////      x63y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9106_1 ( .OUT(na9106_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9106_6 ( .RAM_O1(na9106_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9106_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9107_4 ( .OUT(na9107_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9107_6 ( .RAM_O2(na9107_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9107_2), .COMP_OUT(1'b0) );
// C_AND////      x61y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9108_1 ( .OUT(na9108_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9108_6 ( .RAM_O1(na9108_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9108_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x61y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9109_4 ( .OUT(na9109_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9109_6 ( .RAM_O2(na9109_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9109_2), .COMP_OUT(1'b0) );
// C_AND////      x61y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9110_1 ( .OUT(na9110_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9110_6 ( .RAM_O1(na9110_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9110_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9111_4 ( .OUT(na9111_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9111_6 ( .RAM_O2(na9111_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9111_2), .COMP_OUT(1'b0) );
// C_AND////      x63y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9112_1 ( .OUT(na9112_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9112_6 ( .RAM_O1(na9112_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9112_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9113_4 ( .OUT(na9113_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9113_6 ( .RAM_O2(na9113_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9113_2), .COMP_OUT(1'b0) );
// C_AND////      x63y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9114_1 ( .OUT(na9114_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9114_6 ( .RAM_O1(na9114_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9114_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x63y54     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9115_4 ( .OUT(na9115_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9115_6 ( .RAM_O2(na9115_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na9115_2), .COMP_OUT(1'b0) );
// C_AND////      x63y54     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9116_1 ( .OUT(na9116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a9116_6 ( .RAM_O1(na9116_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na9116_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_////RAM_I2      x66y60     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9117_5 ( .OUT(na9117_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_93), .CP_O(1'b0) );
// C_/RAM_I1///      x66y60     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9118_2 ( .OUT(na9118_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_94), .CP_O(1'b0) );
// C_////RAM_I2      x66y59     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9119_5 ( .OUT(na9119_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_95), .CP_O(1'b0) );
// C_/RAM_I1///      x66y59     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9120_2 ( .OUT(na9120_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_96), .CP_O(1'b0) );
// C_////RAM_I2      x66y58     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9121_5 ( .OUT(na9121_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_97), .CP_O(1'b0) );
// C_/RAM_I1///      x66y58     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9122_2 ( .OUT(na9122_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_98), .CP_O(1'b0) );
// C_////RAM_I2      x66y57     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9123_5 ( .OUT(na9123_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_99), .CP_O(1'b0) );
// C_/RAM_I1///      x66y57     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9124_2 ( .OUT(na9124_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_100), .CP_O(1'b0) );
// C_////RAM_I2      x66y52     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9125_5 ( .OUT(na9125_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_113), .CP_O(1'b0) );
// C_/RAM_I1///      x66y52     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9126_2 ( .OUT(na9126_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_114), .CP_O(1'b0) );
// C_////RAM_I2      x66y51     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9127_5 ( .OUT(na9127_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_115), .CP_O(1'b0) );
// C_/RAM_I1///      x66y51     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9128_2 ( .OUT(na9128_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_116), .CP_O(1'b0) );
// C_////RAM_I2      x66y50     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9129_5 ( .OUT(na9129_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_117), .CP_O(1'b0) );
// C_/RAM_I1///      x66y50     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9130_2 ( .OUT(na9130_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_118), .CP_O(1'b0) );
// C_////RAM_I2      x66y49     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9131_5 ( .OUT(na9131_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_119), .CP_O(1'b0) );
// C_/RAM_I1///      x66y49     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a9132_2 ( .OUT(na9132_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na6659_120), .CP_O(1'b0) );
// C_////Bridge      x111y103     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9133_5 ( .OUT(na9133_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8_2), .IN8(1'b0) );
// C_////Bridge      x90y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9134_5 ( .OUT(na9134_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na9_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y84     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9135_5 ( .OUT(na9135_2), .IN1(1'b0), .IN2(na12_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y71     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9136_5 ( .OUT(na9136_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na18_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9137_5 ( .OUT(na9137_2), .IN1(na19_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y82     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9138_5 ( .OUT(na9138_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na22_1), .IN8(1'b0) );
// C_////Bridge      x81y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9139_5 ( .OUT(na9139_2), .IN1(1'b0), .IN2(na25_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9140_5 ( .OUT(na9140_2), .IN1(1'b0), .IN2(na27_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y78     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9141_5 ( .OUT(na9141_2), .IN1(1'b0), .IN2(na27_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y70     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9142_5 ( .OUT(na9142_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na30_1), .IN8(1'b0) );
// C_////Bridge      x75y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9143_5 ( .OUT(na9143_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na34_2), .IN8(1'b0) );
// C_////Bridge      x88y69     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9144_5 ( .OUT(na9144_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na35_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y65     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9145_5 ( .OUT(na9145_2), .IN1(1'b0), .IN2(na36_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9146_5 ( .OUT(na9146_2), .IN1(1'b0), .IN2(na36_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9147_5 ( .OUT(na9147_2), .IN1(1'b0), .IN2(na36_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9148_5 ( .OUT(na9148_2), .IN1(1'b0), .IN2(na36_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y68     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9149_5 ( .OUT(na9149_2), .IN1(1'b0), .IN2(na36_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y62     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9150_5 ( .OUT(na9150_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na37_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9151_5 ( .OUT(na9151_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na42_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y68     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9152_5 ( .OUT(na9152_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na50_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y70     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9153_5 ( .OUT(na9153_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na61_1) );
// C_////Bridge      x89y74     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9154_5 ( .OUT(na9154_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na66_1), .IN8(1'b0) );
// C_////Bridge      x102y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9155_5 ( .OUT(na9155_2), .IN1(1'b0), .IN2(na67_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9156_5 ( .OUT(na9156_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na73_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9157_5 ( .OUT(na9157_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na73_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9158_5 ( .OUT(na9158_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na73_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y63     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9159_5 ( .OUT(na9159_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na82_1), .IN8(1'b0) );
// C_////Bridge      x84y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9160_5 ( .OUT(na9160_2), .IN1(na86_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y82     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9161_5 ( .OUT(na9161_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na87_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y66     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9162_5 ( .OUT(na9162_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na89_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y56     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9163_5 ( .OUT(na9163_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na89_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y85     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9164_5 ( .OUT(na9164_2), .IN1(1'b0), .IN2(1'b0), .IN3(na90_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9165_5 ( .OUT(na9165_2), .IN1(1'b0), .IN2(1'b0), .IN3(na90_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9166_5 ( .OUT(na9166_2), .IN1(1'b0), .IN2(1'b0), .IN3(na90_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9167_5 ( .OUT(na9167_2), .IN1(1'b0), .IN2(1'b0), .IN3(na90_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y104     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9168_5 ( .OUT(na9168_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na92_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y78     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9169_5 ( .OUT(na9169_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na92_2) );
// C_////Bridge      x90y79     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9170_5 ( .OUT(na9170_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na95_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9171_5 ( .OUT(na9171_2), .IN1(na95_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9172_5 ( .OUT(na9172_2), .IN1(na95_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y81     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9173_5 ( .OUT(na9173_2), .IN1(1'b0), .IN2(1'b0), .IN3(na97_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9174_5 ( .OUT(na9174_2), .IN1(1'b0), .IN2(1'b0), .IN3(na97_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9175_5 ( .OUT(na9175_2), .IN1(1'b0), .IN2(1'b0), .IN3(na97_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9176_5 ( .OUT(na9176_2), .IN1(1'b0), .IN2(1'b0), .IN3(na97_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9177_5 ( .OUT(na9177_2), .IN1(na103_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y87     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9178_5 ( .OUT(na9178_2), .IN1(1'b0), .IN2(1'b0), .IN3(na106_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y76     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9179_5 ( .OUT(na9179_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na154_2) );
// C_////Bridge      x104y67     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9180_5 ( .OUT(na9180_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na155_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9181_5 ( .OUT(na9181_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na160_1) );
// C_////Bridge      x99y77     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9182_5 ( .OUT(na9182_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na165_1) );
// C_////Bridge      x99y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9183_5 ( .OUT(na9183_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na166_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9184_5 ( .OUT(na9184_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na210_1), .IN8(1'b0) );
// C_////Bridge      x97y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9185_5 ( .OUT(na9185_2), .IN1(na214_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9186_5 ( .OUT(na9186_2), .IN1(na214_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9187_5 ( .OUT(na9187_2), .IN1(1'b0), .IN2(na215_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9188_5 ( .OUT(na9188_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na228_1) );
// C_////Bridge      x106y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9189_5 ( .OUT(na9189_2), .IN1(1'b0), .IN2(na267_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y94     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9190_5 ( .OUT(na9190_2), .IN1(1'b0), .IN2(1'b0), .IN3(na278_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y116     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9191_5 ( .OUT(na9191_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na288_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y115     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9192_5 ( .OUT(na9192_2), .IN1(1'b0), .IN2(1'b0), .IN3(na289_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y116     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9193_5 ( .OUT(na9193_2), .IN1(1'b0), .IN2(na291_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y80     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9194_5 ( .OUT(na9194_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na298_1), .IN8(1'b0) );
// C_////Bridge      x94y118     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9195_5 ( .OUT(na9195_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na308_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x133y117     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9196_5 ( .OUT(na9196_2), .IN1(1'b0), .IN2(na316_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y120     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9197_5 ( .OUT(na9197_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na318_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y118     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9198_5 ( .OUT(na9198_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na318_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y120     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9199_5 ( .OUT(na9199_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na324_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y112     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9200_5 ( .OUT(na9200_2), .IN1(1'b0), .IN2(1'b0), .IN3(na336_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9201_5 ( .OUT(na9201_2), .IN1(1'b0), .IN2(na343_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9202_5 ( .OUT(na9202_2), .IN1(1'b0), .IN2(1'b0), .IN3(na347_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9203_5 ( .OUT(na9203_2), .IN1(na356_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y83     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9204_5 ( .OUT(na9204_2), .IN1(1'b0), .IN2(1'b0), .IN3(na359_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9205_5 ( .OUT(na9205_2), .IN1(1'b0), .IN2(1'b0), .IN3(na359_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9206_5 ( .OUT(na9206_2), .IN1(1'b0), .IN2(na369_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y49     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9207_5 ( .OUT(na9207_2), .IN1(1'b0), .IN2(na369_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y91     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9208_5 ( .OUT(na9208_2), .IN1(na374_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9209_5 ( .OUT(na9209_2), .IN1(na374_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y68     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9210_5 ( .OUT(na9210_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na393_2) );
// C_////Bridge      x80y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9211_5 ( .OUT(na9211_2), .IN1(1'b0), .IN2(na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9212_5 ( .OUT(na9212_2), .IN1(1'b0), .IN2(na401_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9213_5 ( .OUT(na9213_2), .IN1(na402_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9214_5 ( .OUT(na9214_2), .IN1(1'b0), .IN2(1'b0), .IN3(na403_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9215_5 ( .OUT(na9215_2), .IN1(1'b0), .IN2(1'b0), .IN3(na403_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y99     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9216_5 ( .OUT(na9216_2), .IN1(1'b0), .IN2(1'b0), .IN3(na403_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9217_5 ( .OUT(na9217_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na406_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9218_5 ( .OUT(na9218_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na406_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9219_5 ( .OUT(na9219_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na406_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y99     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9220_5 ( .OUT(na9220_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na410_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y60     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9221_5 ( .OUT(na9221_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na423_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y81     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9222_5 ( .OUT(na9222_2), .IN1(na428_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9223_5 ( .OUT(na9223_2), .IN1(na428_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9224_5 ( .OUT(na9224_2), .IN1(na428_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y78     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9225_5 ( .OUT(na9225_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na432_1), .IN8(1'b0) );
// C_////Bridge      x91y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9226_5 ( .OUT(na9226_2), .IN1(1'b0), .IN2(na435_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9227_5 ( .OUT(na9227_2), .IN1(1'b0), .IN2(na435_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y84     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9228_5 ( .OUT(na9228_2), .IN1(1'b0), .IN2(na435_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9229_5 ( .OUT(na9229_2), .IN1(1'b0), .IN2(1'b0), .IN3(na436_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9230_5 ( .OUT(na9230_2), .IN1(1'b0), .IN2(1'b0), .IN3(na436_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y89     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9231_5 ( .OUT(na9231_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na452_1) );
// C_////Bridge      x93y87     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9232_5 ( .OUT(na9232_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na452_2) );
// C_////Bridge      x92y74     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9233_5 ( .OUT(na9233_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na456_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9234_5 ( .OUT(na9234_2), .IN1(na457_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y77     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9235_5 ( .OUT(na9235_2), .IN1(1'b0), .IN2(na459_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y93     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9236_5 ( .OUT(na9236_2), .IN1(na463_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y75     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9237_5 ( .OUT(na9237_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na478_2), .IN8(1'b0) );
// C_////Bridge      x104y88     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9238_5 ( .OUT(na9238_2), .IN1(1'b0), .IN2(na483_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9239_5 ( .OUT(na9239_2), .IN1(1'b0), .IN2(na486_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9240_5 ( .OUT(na9240_2), .IN1(1'b0), .IN2(na486_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9241_5 ( .OUT(na9241_2), .IN1(na488_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9242_5 ( .OUT(na9242_2), .IN1(na488_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y64     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9243_5 ( .OUT(na9243_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na488_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9244_5 ( .OUT(na9244_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na500_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9245_5 ( .OUT(na9245_2), .IN1(1'b0), .IN2(na504_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9246_5 ( .OUT(na9246_2), .IN1(1'b0), .IN2(1'b0), .IN3(na517_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9247_5 ( .OUT(na9247_2), .IN1(1'b0), .IN2(1'b0), .IN3(na517_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9248_5 ( .OUT(na9248_2), .IN1(1'b0), .IN2(1'b0), .IN3(na517_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9249_5 ( .OUT(na9249_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na523_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9250_5 ( .OUT(na9250_2), .IN1(na528_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9251_5 ( .OUT(na9251_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na533_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y108     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9252_5 ( .OUT(na9252_2), .IN1(1'b0), .IN2(na536_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y61     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9253_5 ( .OUT(na9253_2), .IN1(na540_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9254_5 ( .OUT(na9254_2), .IN1(na540_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y122     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9255_5 ( .OUT(na9255_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na542_1), .IN8(1'b0) );
// C_////Bridge      x53y65     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9256_5 ( .OUT(na9256_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na545_1), .IN8(1'b0) );
// C_////Bridge      x68y122     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9257_5 ( .OUT(na9257_2), .IN1(na546_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9258_5 ( .OUT(na9258_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na546_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y108     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9259_5 ( .OUT(na9259_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na547_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9260_5 ( .OUT(na9260_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na547_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9261_5 ( .OUT(na9261_2), .IN1(1'b0), .IN2(1'b0), .IN3(na550_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y108     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9262_5 ( .OUT(na9262_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na552_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9263_5 ( .OUT(na9263_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na552_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9264_5 ( .OUT(na9264_2), .IN1(1'b0), .IN2(1'b0), .IN3(na561_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9265_5 ( .OUT(na9265_2), .IN1(na566_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y79     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9266_5 ( .OUT(na9266_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na567_1), .IN8(1'b0) );
// C_////Bridge      x112y84     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9267_5 ( .OUT(na9267_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na570_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9268_5 ( .OUT(na9268_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na574_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9269_5 ( .OUT(na9269_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na574_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y84     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9270_5 ( .OUT(na9270_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na579_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y123     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9271_5 ( .OUT(na9271_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na587_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9272_5 ( .OUT(na9272_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na588_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y121     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9273_5 ( .OUT(na9273_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na588_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y62     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9274_5 ( .OUT(na9274_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na589_1), .IN8(1'b0) );
// C_////Bridge      x51y59     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9275_5 ( .OUT(na9275_2), .IN1(1'b0), .IN2(1'b0), .IN3(na589_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9276_5 ( .OUT(na9276_2), .IN1(na590_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9277_5 ( .OUT(na9277_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na597_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y116     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9278_5 ( .OUT(na9278_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na598_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y123     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9279_5 ( .OUT(na9279_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na598_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9280_5 ( .OUT(na9280_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na603_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9281_5 ( .OUT(na9281_2), .IN1(1'b0), .IN2(1'b0), .IN3(na607_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9282_5 ( .OUT(na9282_2), .IN1(1'b0), .IN2(1'b0), .IN3(na608_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y121     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9283_5 ( .OUT(na9283_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na609_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y110     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9284_5 ( .OUT(na9284_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na614_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9285_5 ( .OUT(na9285_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na614_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y66     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9286_5 ( .OUT(na9286_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na617_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y118     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9287_5 ( .OUT(na9287_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na619_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y121     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9288_5 ( .OUT(na9288_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na619_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y106     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9289_5 ( .OUT(na9289_2), .IN1(na620_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9290_5 ( .OUT(na9290_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na624_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9291_5 ( .OUT(na9291_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na624_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9292_5 ( .OUT(na9292_2), .IN1(1'b0), .IN2(1'b0), .IN3(na632_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9293_5 ( .OUT(na9293_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na633_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y112     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9294_5 ( .OUT(na9294_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na634_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y123     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9295_5 ( .OUT(na9295_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na634_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9296_5 ( .OUT(na9296_2), .IN1(na643_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y88     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9297_5 ( .OUT(na9297_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na652_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y93     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9298_5 ( .OUT(na9298_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na654_1) );
// C_////Bridge      x55y112     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9299_5 ( .OUT(na9299_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na658_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9300_5 ( .OUT(na9300_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na658_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y81     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9301_5 ( .OUT(na9301_2), .IN1(1'b0), .IN2(1'b0), .IN3(na661_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y85     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9302_5 ( .OUT(na9302_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na663_1) );
// C_////Bridge      x57y116     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9303_5 ( .OUT(na9303_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na664_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9304_5 ( .OUT(na9304_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na664_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y121     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9305_5 ( .OUT(na9305_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na673_2) );
// C_////Bridge      x64y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9306_5 ( .OUT(na9306_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na678_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y112     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9307_5 ( .OUT(na9307_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na679_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y123     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9308_5 ( .OUT(na9308_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na679_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y121     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9309_5 ( .OUT(na9309_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na684_1) );
// C_////Bridge      x58y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9310_5 ( .OUT(na9310_2), .IN1(na687_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9311_5 ( .OUT(na9311_2), .IN1(na687_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y123     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9312_5 ( .OUT(na9312_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na689_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y122     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9313_5 ( .OUT(na9313_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na694_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9314_5 ( .OUT(na9314_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na694_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y73     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9315_5 ( .OUT(na9315_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na697_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y116     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9316_5 ( .OUT(na9316_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na699_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9317_5 ( .OUT(na9317_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na699_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9318_5 ( .OUT(na9318_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na707_1), .IN8(1'b0) );
// C_////Bridge      x68y117     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9319_5 ( .OUT(na9319_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na708_2) );
// C_////Bridge      x73y96     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9320_5 ( .OUT(na9320_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na714_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y116     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9321_5 ( .OUT(na9321_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na719_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y121     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9322_5 ( .OUT(na9322_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na719_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y62     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9323_5 ( .OUT(na9323_2), .IN1(1'b0), .IN2(na728_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y93     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9324_5 ( .OUT(na9324_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na731_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y110     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9325_5 ( .OUT(na9325_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na731_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y64     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9326_5 ( .OUT(na9326_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na737_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y61     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9327_5 ( .OUT(na9327_2), .IN1(na745_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x135y101     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9328_5 ( .OUT(na9328_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na755_2), .IN8(1'b0) );
// C_////Bridge      x93y95     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9329_5 ( .OUT(na9329_2), .IN1(1'b0), .IN2(1'b0), .IN3(na757_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y84     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9330_5 ( .OUT(na9330_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na758_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y66     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9331_5 ( .OUT(na9331_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na767_2) );
// C_////Bridge      x79y66     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9332_5 ( .OUT(na9332_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na771_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y64     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9333_5 ( .OUT(na9333_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na775_2) );
// C_////Bridge      x111y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9334_5 ( .OUT(na9334_2), .IN1(1'b0), .IN2(na785_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y83     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9335_5 ( .OUT(na9335_2), .IN1(1'b0), .IN2(1'b0), .IN3(na791_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9336_5 ( .OUT(na9336_2), .IN1(1'b0), .IN2(1'b0), .IN3(na791_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y76     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9337_5 ( .OUT(na9337_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na798_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y93     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9338_5 ( .OUT(na9338_2), .IN1(na799_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y99     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9339_5 ( .OUT(na9339_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na803_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y81     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9340_5 ( .OUT(na9340_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na827_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9341_5 ( .OUT(na9341_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na834_2) );
// C_////Bridge      x88y72     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9342_5 ( .OUT(na9342_2), .IN1(1'b0), .IN2(na843_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y80     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9343_5 ( .OUT(na9343_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na847_2) );
// C_////Bridge      x98y107     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9344_5 ( .OUT(na9344_2), .IN1(na853_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y110     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9345_5 ( .OUT(na9345_2), .IN1(na853_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y75     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9346_5 ( .OUT(na9346_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na857_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y82     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9347_5 ( .OUT(na9347_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na870_1) );
// C_////Bridge      x77y82     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9348_5 ( .OUT(na9348_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na870_2) );
// C_////Bridge      x107y83     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9349_5 ( .OUT(na9349_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na892_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y105     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9350_5 ( .OUT(na9350_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na894_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9351_5 ( .OUT(na9351_2), .IN1(1'b0), .IN2(1'b0), .IN3(na903_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9352_5 ( .OUT(na9352_2), .IN1(na906_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y106     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9353_5 ( .OUT(na9353_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na913_1), .IN8(1'b0) );
// C_////Bridge      x93y107     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9354_5 ( .OUT(na9354_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na913_2), .IN8(1'b0) );
// C_////Bridge      x92y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9355_5 ( .OUT(na9355_2), .IN1(1'b0), .IN2(na916_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y104     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9356_5 ( .OUT(na9356_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na925_1), .IN8(1'b0) );
// C_////Bridge      x91y105     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9357_5 ( .OUT(na9357_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na925_2), .IN8(1'b0) );
// C_////Bridge      x104y92     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9358_5 ( .OUT(na9358_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na936_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y70     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9359_5 ( .OUT(na9359_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na947_1) );
// C_////Bridge      x89y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9360_5 ( .OUT(na9360_2), .IN1(1'b0), .IN2(na955_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9361_5 ( .OUT(na9361_2), .IN1(1'b0), .IN2(na955_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9362_5 ( .OUT(na9362_2), .IN1(1'b0), .IN2(na955_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y68     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9363_5 ( .OUT(na9363_2), .IN1(1'b0), .IN2(na958_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9364_5 ( .OUT(na9364_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na973_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y56     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9365_5 ( .OUT(na9365_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na973_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9366_5 ( .OUT(na9366_2), .IN1(1'b0), .IN2(1'b0), .IN3(na977_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y59     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9367_5 ( .OUT(na9367_2), .IN1(1'b0), .IN2(1'b0), .IN3(na977_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9368_5 ( .OUT(na9368_2), .IN1(1'b0), .IN2(1'b0), .IN3(na977_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9369_5 ( .OUT(na9369_2), .IN1(1'b0), .IN2(na980_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9370_5 ( .OUT(na9370_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na981_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y45     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9371_5 ( .OUT(na9371_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na985_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x131y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9372_5 ( .OUT(na9372_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na989_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9373_5 ( .OUT(na9373_2), .IN1(1'b0), .IN2(1'b0), .IN3(na997_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y90     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9374_5 ( .OUT(na9374_2), .IN1(1'b0), .IN2(1'b0), .IN3(na997_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y74     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9375_5 ( .OUT(na9375_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1001_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y84     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9376_5 ( .OUT(na9376_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1010_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9377_5 ( .OUT(na9377_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1016_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y101     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9378_5 ( .OUT(na9378_2), .IN1(na1022_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y110     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9379_5 ( .OUT(na9379_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1033_1), .IN8(1'b0) );
// C_////Bridge      x112y106     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9380_5 ( .OUT(na9380_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1035_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y89     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9381_5 ( .OUT(na9381_2), .IN1(na1039_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y85     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9382_5 ( .OUT(na9382_2), .IN1(na1045_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9383_5 ( .OUT(na9383_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1054_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y72     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9384_5 ( .OUT(na9384_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1054_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y104     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9385_5 ( .OUT(na9385_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1061_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y103     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9386_5 ( .OUT(na9386_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1061_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y97     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9387_5 ( .OUT(na9387_2), .IN1(1'b0), .IN2(na1064_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9388_5 ( .OUT(na9388_2), .IN1(1'b0), .IN2(na1064_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y104     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9389_5 ( .OUT(na9389_2), .IN1(1'b0), .IN2(na1064_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y88     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9390_5 ( .OUT(na9390_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1065_1), .IN8(1'b0) );
// C_////Bridge      x89y83     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9391_5 ( .OUT(na9391_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1065_2), .IN8(1'b0) );
// C_////Bridge      x114y108     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9392_5 ( .OUT(na9392_2), .IN1(na1069_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y110     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9393_5 ( .OUT(na9393_2), .IN1(na1070_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y107     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9394_5 ( .OUT(na9394_2), .IN1(1'b0), .IN2(na1074_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y82     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9395_5 ( .OUT(na9395_2), .IN1(na1076_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y84     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9396_5 ( .OUT(na9396_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1079_1) );
// C_////Bridge      x110y94     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9397_5 ( .OUT(na9397_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1081_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9398_5 ( .OUT(na9398_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1085_1), .IN8(1'b0) );
// C_////Bridge      x122y110     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9399_5 ( .OUT(na9399_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1087_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y101     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9400_5 ( .OUT(na9400_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1088_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y108     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9401_5 ( .OUT(na9401_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1088_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y106     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9402_5 ( .OUT(na9402_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1094_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y99     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9403_5 ( .OUT(na9403_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1096_1), .IN8(1'b0) );
// C_////Bridge      x99y90     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9404_5 ( .OUT(na9404_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1113_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9405_5 ( .OUT(na9405_2), .IN1(na1115_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y106     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9406_5 ( .OUT(na9406_2), .IN1(na1115_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y102     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9407_5 ( .OUT(na9407_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1117_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y95     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9408_5 ( .OUT(na9408_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1118_1), .IN8(1'b0) );
// C_////Bridge      x123y105     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9409_5 ( .OUT(na9409_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1121_1) );
// C_////Bridge      x120y96     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9410_5 ( .OUT(na9410_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1123_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y60     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9411_5 ( .OUT(na9411_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1130_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9412_5 ( .OUT(na9412_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1134_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9413_5 ( .OUT(na9413_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1135_1) );
// C_////Bridge      x99y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9414_5 ( .OUT(na9414_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1136_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9415_5 ( .OUT(na9415_2), .IN1(na1138_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y100     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9416_5 ( .OUT(na9416_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1145_1), .IN8(1'b0) );
// C_////Bridge      x109y107     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9417_5 ( .OUT(na9417_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1147_1) );
// C_////Bridge      x106y99     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9418_5 ( .OUT(na9418_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1149_1) );
// C_////Bridge      x113y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9419_5 ( .OUT(na9419_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1150_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9420_5 ( .OUT(na9420_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1150_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y105     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9421_5 ( .OUT(na9421_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1153_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y98     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9422_5 ( .OUT(na9422_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1153_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9423_5 ( .OUT(na9423_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1154_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y106     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9424_5 ( .OUT(na9424_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1154_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y94     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9425_5 ( .OUT(na9425_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1155_1) );
// C_////Bridge      x103y91     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9426_5 ( .OUT(na9426_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1156_1) );
// C_////Bridge      x95y97     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9427_5 ( .OUT(na9427_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1157_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9428_5 ( .OUT(na9428_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1157_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y93     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9429_5 ( .OUT(na9429_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1158_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y104     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9430_5 ( .OUT(na9430_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1158_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9431_5 ( .OUT(na9431_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1159_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9432_5 ( .OUT(na9432_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1162_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y109     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9433_5 ( .OUT(na9433_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1162_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y107     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9434_5 ( .OUT(na9434_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1163_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y110     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9435_5 ( .OUT(na9435_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1164_1) );
// C_////Bridge      x102y59     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9436_5 ( .OUT(na9436_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1171_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y61     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9437_5 ( .OUT(na9437_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1172_1) );
// C_////Bridge      x93y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9438_5 ( .OUT(na9438_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1175_1) );
// C_////Bridge      x71y86     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9439_5 ( .OUT(na9439_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1175_2) );
// C_////Bridge      x86y92     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9440_5 ( .OUT(na9440_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1177_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y95     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9441_5 ( .OUT(na9441_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1181_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9442_5 ( .OUT(na9442_2), .IN1(na1187_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y113     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9443_5 ( .OUT(na9443_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1197_1) );
// C_////Bridge      x107y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9444_5 ( .OUT(na9444_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1198_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9445_5 ( .OUT(na9445_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1198_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y109     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9446_5 ( .OUT(na9446_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1199_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9447_5 ( .OUT(na9447_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1199_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y107     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9448_5 ( .OUT(na9448_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1200_1) );
// C_////Bridge      x108y100     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9449_5 ( .OUT(na9449_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1202_1), .IN8(1'b0) );
// C_////Bridge      x105y107     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9450_5 ( .OUT(na9450_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1203_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y107     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9451_5 ( .OUT(na9451_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1203_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y111     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9452_5 ( .OUT(na9452_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1204_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y112     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9453_5 ( .OUT(na9453_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1205_1) );
// C_////Bridge      x99y109     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9454_5 ( .OUT(na9454_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1206_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9455_5 ( .OUT(na9455_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1206_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y111     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9456_5 ( .OUT(na9456_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1207_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y107     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9457_5 ( .OUT(na9457_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1207_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y111     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9458_5 ( .OUT(na9458_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1208_1) );
// C_////Bridge      x105y113     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9459_5 ( .OUT(na9459_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1209_1) );
// C_////Bridge      x113y111     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9460_5 ( .OUT(na9460_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1210_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y103     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9461_5 ( .OUT(na9461_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1210_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9462_5 ( .OUT(na9462_2), .IN1(na1222_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9463_5 ( .OUT(na9463_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1223_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y91     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9464_5 ( .OUT(na9464_2), .IN1(na1225_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y115     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9465_5 ( .OUT(na9465_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1227_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y112     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9466_5 ( .OUT(na9466_2), .IN1(1'b0), .IN2(na1228_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y113     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9467_5 ( .OUT(na9467_2), .IN1(1'b0), .IN2(na1229_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9468_5 ( .OUT(na9468_2), .IN1(1'b0), .IN2(na1232_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y121     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9469_5 ( .OUT(na9469_2), .IN1(1'b0), .IN2(na1233_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y120     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9470_5 ( .OUT(na9470_2), .IN1(1'b0), .IN2(na1234_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y119     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9471_5 ( .OUT(na9471_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1238_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y119     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9472_5 ( .OUT(na9472_2), .IN1(1'b0), .IN2(na1241_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y120     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9473_5 ( .OUT(na9473_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1242_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y111     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9474_5 ( .OUT(na9474_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1243_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y113     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9475_5 ( .OUT(na9475_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1245_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9476_5 ( .OUT(na9476_2), .IN1(na1246_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y117     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9477_5 ( .OUT(na9477_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1261_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y116     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9478_5 ( .OUT(na9478_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1262_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9479_5 ( .OUT(na9479_2), .IN1(1'b0), .IN2(na1263_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y100     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9480_5 ( .OUT(na9480_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1265_1) );
// C_////Bridge      x110y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9481_5 ( .OUT(na9481_2), .IN1(1'b0), .IN2(na1266_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y92     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9482_5 ( .OUT(na9482_2), .IN1(1'b0), .IN2(na1267_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9483_5 ( .OUT(na9483_2), .IN1(1'b0), .IN2(na1268_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y115     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9484_5 ( .OUT(na9484_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1269_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y118     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9485_5 ( .OUT(na9485_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1272_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y104     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9486_5 ( .OUT(na9486_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1314_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y101     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9487_5 ( .OUT(na9487_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1314_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9488_5 ( .OUT(na9488_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1337_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y101     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9489_5 ( .OUT(na9489_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1337_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y82     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9490_5 ( .OUT(na9490_2), .IN1(na1342_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y97     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9491_5 ( .OUT(na9491_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1346_1) );
// C_////Bridge      x94y85     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9492_5 ( .OUT(na9492_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1351_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y85     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9493_5 ( .OUT(na9493_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1353_1) );
// C_////Bridge      x110y104     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9494_5 ( .OUT(na9494_2), .IN1(na1354_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9495_5 ( .OUT(na9495_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1355_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y77     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9496_5 ( .OUT(na9496_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1355_2), .IN8(1'b0) );
// C_////Bridge      x87y86     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9497_5 ( .OUT(na9497_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1359_1), .IN8(1'b0) );
// C_////Bridge      x91y83     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9498_5 ( .OUT(na9498_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1359_2), .IN8(1'b0) );
// C_////Bridge      x115y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9499_5 ( .OUT(na9499_2), .IN1(1'b0), .IN2(na1371_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9500_5 ( .OUT(na9500_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1377_1) );
// C_////Bridge      x113y89     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9501_5 ( .OUT(na9501_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1382_1) );
// C_////Bridge      x65y64     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9502_5 ( .OUT(na9502_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1387_2), .IN8(1'b0) );
// C_////Bridge      x69y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9503_5 ( .OUT(na9503_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1407_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9504_5 ( .OUT(na9504_2), .IN1(1'b0), .IN2(na1411_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y81     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9505_5 ( .OUT(na9505_2), .IN1(na1416_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y42     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9506_5 ( .OUT(na9506_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1425_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y37     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9507_5 ( .OUT(na9507_2), .IN1(na1427_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y41     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9508_5 ( .OUT(na9508_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1427_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y96     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9509_5 ( .OUT(na9509_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1433_1), .IN8(1'b0) );
// C_////Bridge      x116y71     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9510_5 ( .OUT(na9510_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1447_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9511_5 ( .OUT(na9511_2), .IN1(1'b0), .IN2(na1462_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y92     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9512_5 ( .OUT(na9512_2), .IN1(1'b0), .IN2(na1462_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y94     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9513_5 ( .OUT(na9513_2), .IN1(1'b0), .IN2(na1462_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y92     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9514_5 ( .OUT(na9514_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1481_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y76     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9515_5 ( .OUT(na9515_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1498_2), .IN8(1'b0) );
// C_////Bridge      x123y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9516_5 ( .OUT(na9516_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1512_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y87     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9517_5 ( .OUT(na9517_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1512_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y76     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9518_5 ( .OUT(na9518_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1525_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y79     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9519_5 ( .OUT(na9519_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1527_1) );
// C_////Bridge      x55y116     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9520_5 ( .OUT(na9520_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1583_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9521_5 ( .OUT(na9521_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1583_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y73     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9522_5 ( .OUT(na9522_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1586_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9523_5 ( .OUT(na9523_2), .IN1(1'b0), .IN2(na1595_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y108     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9524_5 ( .OUT(na9524_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1600_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9525_5 ( .OUT(na9525_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1600_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y67     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9526_5 ( .OUT(na9526_2), .IN1(na1603_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y75     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9527_5 ( .OUT(na9527_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1623_1) );
// C_////Bridge      x98y100     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9528_5 ( .OUT(na9528_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1656_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9529_5 ( .OUT(na9529_2), .IN1(na1658_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9530_5 ( .OUT(na9530_2), .IN1(1'b0), .IN2(na1693_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y103     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9531_5 ( .OUT(na9531_2), .IN1(na1695_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y88     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9532_5 ( .OUT(na9532_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1726_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y65     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9533_5 ( .OUT(na9533_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1770_2) );
// C_////Bridge      x91y61     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9534_5 ( .OUT(na9534_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1858_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y42     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9535_5 ( .OUT(na9535_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1865_1) );
// C_////Bridge      x104y71     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9536_5 ( .OUT(na9536_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1885_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9537_5 ( .OUT(na9537_2), .IN1(na1889_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9538_5 ( .OUT(na9538_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1891_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9539_5 ( .OUT(na9539_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1894_1) );
// C_////Bridge      x100y100     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9540_5 ( .OUT(na9540_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1903_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y65     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9541_5 ( .OUT(na9541_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1921_1) );
// C_////Bridge      x89y72     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9542_5 ( .OUT(na9542_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1921_2) );
// C_////Bridge      x86y43     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9543_5 ( .OUT(na9543_2), .IN1(na1960_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y60     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9544_5 ( .OUT(na9544_2), .IN1(na1978_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y56     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9545_5 ( .OUT(na9545_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1987_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9546_5 ( .OUT(na9546_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1994_2) );
// C_////Bridge      x83y38     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9547_5 ( .OUT(na9547_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2001_2) );
// C_////Bridge      x84y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9548_5 ( .OUT(na9548_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2004_1) );
// C_////Bridge      x87y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9549_5 ( .OUT(na9549_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2015_2) );
// C_////Bridge      x87y44     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9550_5 ( .OUT(na9550_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2022_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y44     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9551_5 ( .OUT(na9551_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2029_2) );
// C_////Bridge      x86y59     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9552_5 ( .OUT(na9552_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2036_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9553_5 ( .OUT(na9553_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2064_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y72     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9554_5 ( .OUT(na9554_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2078_2) );
// C_////Bridge      x85y60     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9555_5 ( .OUT(na9555_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2099_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y38     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9556_5 ( .OUT(na9556_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2106_2) );
// C_////Bridge      x87y38     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9557_5 ( .OUT(na9557_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2113_2) );
// C_////Bridge      x85y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9558_5 ( .OUT(na9558_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2120_2) );
// C_////Bridge      x89y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9559_5 ( .OUT(na9559_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2127_2) );
// C_////Bridge      x87y42     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9560_5 ( .OUT(na9560_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2134_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9561_5 ( .OUT(na9561_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2136_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y42     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9562_5 ( .OUT(na9562_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2141_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9563_5 ( .OUT(na9563_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2143_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y79     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9564_5 ( .OUT(na9564_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2168_1) );
// C_////Bridge      x65y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9565_5 ( .OUT(na9565_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2171_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y119     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9566_5 ( .OUT(na9566_2), .IN1(1'b0), .IN2(na2172_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9567_5 ( .OUT(na9567_2), .IN1(na2246_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y69     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9568_5 ( .OUT(na9568_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2309_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9569_5 ( .OUT(na9569_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2311_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9570_5 ( .OUT(na9570_2), .IN1(1'b0), .IN2(na2314_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9571_5 ( .OUT(na9571_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2316_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9572_5 ( .OUT(na9572_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2316_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9573_5 ( .OUT(na9573_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2318_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9574_5 ( .OUT(na9574_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2321_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9575_5 ( .OUT(na9575_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2327_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9576_5 ( .OUT(na9576_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2327_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9577_5 ( .OUT(na9577_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2327_2), .IN8(1'b0) );
// C_////Bridge      x50y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9578_5 ( .OUT(na9578_2), .IN1(na2332_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9579_5 ( .OUT(na9579_2), .IN1(na2332_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y63     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9580_5 ( .OUT(na9580_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2335_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9581_5 ( .OUT(na9581_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2335_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9582_5 ( .OUT(na9582_2), .IN1(1'b0), .IN2(na2340_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y59     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9583_5 ( .OUT(na9583_2), .IN1(1'b0), .IN2(na2340_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y75     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9584_5 ( .OUT(na9584_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2348_1) );
// C_////Bridge      x51y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9585_5 ( .OUT(na9585_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2357_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y69     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9586_5 ( .OUT(na9586_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2357_2), .IN8(1'b0) );
// C_////Bridge      x57y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9587_5 ( .OUT(na9587_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2369_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9588_5 ( .OUT(na9588_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2369_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9589_5 ( .OUT(na9589_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2369_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9590_5 ( .OUT(na9590_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2372_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y74     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9591_5 ( .OUT(na9591_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2372_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y61     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9592_5 ( .OUT(na9592_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2372_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9593_5 ( .OUT(na9593_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2372_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y78     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9594_5 ( .OUT(na9594_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2390_1), .IN8(1'b0) );
// C_////Bridge      x68y82     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9595_5 ( .OUT(na9595_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2391_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9596_5 ( .OUT(na9596_2), .IN1(na2392_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9597_5 ( .OUT(na9597_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2395_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9598_5 ( .OUT(na9598_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2398_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9599_5 ( .OUT(na9599_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2400_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y86     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9600_5 ( .OUT(na9600_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2407_1), .IN8(1'b0) );
// C_////Bridge      x59y87     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9601_5 ( .OUT(na9601_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2408_1), .IN8(1'b0) );
// C_////Bridge      x57y94     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9602_5 ( .OUT(na9602_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2419_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y78     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9603_5 ( .OUT(na9603_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2422_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y62     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9604_5 ( .OUT(na9604_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2425_2) );
// C_////Bridge      x73y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9605_5 ( .OUT(na9605_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2427_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9606_5 ( .OUT(na9606_2), .IN1(1'b0), .IN2(na2429_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y65     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9607_5 ( .OUT(na9607_2), .IN1(1'b0), .IN2(na2433_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y67     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9608_5 ( .OUT(na9608_2), .IN1(1'b0), .IN2(na2434_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y89     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9609_5 ( .OUT(na9609_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2440_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9610_5 ( .OUT(na9610_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2441_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y90     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9611_5 ( .OUT(na9611_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2442_1), .IN8(1'b0) );
// C_////Bridge      x58y90     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9612_5 ( .OUT(na9612_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2443_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y59     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9613_5 ( .OUT(na9613_2), .IN1(1'b0), .IN2(na2457_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y80     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9614_5 ( .OUT(na9614_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2555_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y74     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9615_5 ( .OUT(na9615_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2556_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9616_5 ( .OUT(na9616_2), .IN1(1'b0), .IN2(na2557_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9617_5 ( .OUT(na9617_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2558_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9618_5 ( .OUT(na9618_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2558_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9619_5 ( .OUT(na9619_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2558_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9620_5 ( .OUT(na9620_2), .IN1(na2562_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9621_5 ( .OUT(na9621_2), .IN1(1'b0), .IN2(na2564_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y79     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9622_5 ( .OUT(na9622_2), .IN1(na2565_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9623_5 ( .OUT(na9623_2), .IN1(na2565_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y98     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9624_5 ( .OUT(na9624_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2568_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y86     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9625_5 ( .OUT(na9625_2), .IN1(1'b0), .IN2(na2571_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9626_5 ( .OUT(na9626_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2572_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y79     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9627_5 ( .OUT(na9627_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2572_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y86     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9628_5 ( .OUT(na9628_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2573_1) );
// C_////Bridge      x75y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9629_5 ( .OUT(na9629_2), .IN1(na2574_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9630_5 ( .OUT(na9630_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2580_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y79     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9631_5 ( .OUT(na9631_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2582_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y86     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9632_5 ( .OUT(na9632_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2594_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y87     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9633_5 ( .OUT(na9633_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2598_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y80     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9634_5 ( .OUT(na9634_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2600_1), .IN8(1'b0) );
// C_////Bridge      x79y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9635_5 ( .OUT(na9635_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2601_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9636_5 ( .OUT(na9636_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2602_1) );
// C_////Bridge      x54y84     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9637_5 ( .OUT(na9637_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2603_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y84     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9638_5 ( .OUT(na9638_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2608_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y89     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9639_5 ( .OUT(na9639_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2609_1) );
// C_////Bridge      x68y70     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9640_5 ( .OUT(na9640_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2610_1), .IN8(1'b0) );
// C_////Bridge      x67y87     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9641_5 ( .OUT(na9641_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2613_1), .IN8(1'b0) );
// C_////Bridge      x59y94     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9642_5 ( .OUT(na9642_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2615_1) );
// C_////Bridge      x57y93     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9643_5 ( .OUT(na9643_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2616_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9644_5 ( .OUT(na9644_2), .IN1(na2622_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y92     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9645_5 ( .OUT(na9645_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2623_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9646_5 ( .OUT(na9646_2), .IN1(1'b0), .IN2(na2626_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y92     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9647_5 ( .OUT(na9647_2), .IN1(1'b0), .IN2(na2626_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y93     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9648_5 ( .OUT(na9648_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2661_1) );
// C_////Bridge      x116y113     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9649_5 ( .OUT(na9649_2), .IN1(1'b0), .IN2(na2666_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9650_5 ( .OUT(na9650_2), .IN1(1'b0), .IN2(na2668_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y104     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9651_5 ( .OUT(na9651_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2670_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y96     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9652_5 ( .OUT(na9652_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2673_1), .IN8(1'b0) );
// C_////Bridge      x91y100     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9653_5 ( .OUT(na9653_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2677_1), .IN8(1'b0) );
// C_////Bridge      x91y99     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9654_5 ( .OUT(na9654_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2677_2), .IN8(1'b0) );
// C_////Bridge      x91y106     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9655_5 ( .OUT(na9655_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2681_1), .IN8(1'b0) );
// C_////Bridge      x93y105     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9656_5 ( .OUT(na9656_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2681_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9657_5 ( .OUT(na9657_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2687_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y81     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9658_5 ( .OUT(na9658_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2687_2), .IN8(1'b0) );
// C_////Bridge      x112y94     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9659_5 ( .OUT(na9659_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2693_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y71     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9660_5 ( .OUT(na9660_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2698_1), .IN8(1'b0) );
// C_////Bridge      x117y99     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9661_5 ( .OUT(na9661_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2701_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y106     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9662_5 ( .OUT(na9662_2), .IN1(na2702_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y86     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9663_5 ( .OUT(na9663_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2703_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y97     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9664_5 ( .OUT(na9664_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2704_1), .IN8(1'b0) );
// C_////Bridge      x132y54     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9665_5 ( .OUT(na9665_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2718_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y105     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9666_5 ( .OUT(na9666_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2721_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y104     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9667_5 ( .OUT(na9667_2), .IN1(na2733_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y95     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9668_5 ( .OUT(na9668_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2740_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9669_5 ( .OUT(na9669_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2740_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9670_5 ( .OUT(na9670_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2750_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y53     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9671_5 ( .OUT(na9671_2), .IN1(1'b0), .IN2(na2759_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y93     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9672_5 ( .OUT(na9672_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2762_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9673_5 ( .OUT(na9673_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2762_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9674_5 ( .OUT(na9674_2), .IN1(1'b0), .IN2(na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9675_5 ( .OUT(na9675_2), .IN1(1'b0), .IN2(na2773_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y69     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9676_5 ( .OUT(na9676_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2781_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9677_5 ( .OUT(na9677_2), .IN1(1'b0), .IN2(na2782_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y70     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9678_5 ( .OUT(na9678_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2783_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y77     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9679_5 ( .OUT(na9679_2), .IN1(1'b0), .IN2(na2784_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y74     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9680_5 ( .OUT(na9680_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2786_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9681_5 ( .OUT(na9681_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2788_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9682_5 ( .OUT(na9682_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2788_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y83     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9683_5 ( .OUT(na9683_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2791_1) );
// C_////Bridge      x107y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9684_5 ( .OUT(na9684_2), .IN1(1'b0), .IN2(na2795_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y79     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9685_5 ( .OUT(na9685_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2798_1) );
// C_////Bridge      x118y82     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9686_5 ( .OUT(na9686_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2802_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y86     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9687_5 ( .OUT(na9687_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2805_1), .IN8(1'b0) );
// C_////Bridge      x109y85     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9688_5 ( .OUT(na9688_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2805_2), .IN8(1'b0) );
// C_////Bridge      x125y96     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9689_5 ( .OUT(na9689_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2811_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y95     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9690_5 ( .OUT(na9690_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2811_2), .IN8(1'b0) );
// C_////Bridge      x107y84     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9691_5 ( .OUT(na9691_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2818_1), .IN8(1'b0) );
// C_////Bridge      x107y81     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9692_5 ( .OUT(na9692_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2818_2), .IN8(1'b0) );
// C_////Bridge      x115y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9693_5 ( .OUT(na9693_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2827_1) );
// C_////Bridge      x110y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9694_5 ( .OUT(na9694_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2829_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9695_5 ( .OUT(na9695_2), .IN1(na2832_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9696_5 ( .OUT(na9696_2), .IN1(1'b0), .IN2(na2834_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y72     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9697_5 ( .OUT(na9697_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2838_1), .IN8(1'b0) );
// C_////Bridge      x53y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9698_5 ( .OUT(na9698_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2840_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9699_5 ( .OUT(na9699_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2845_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y35     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9700_5 ( .OUT(na9700_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2847_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y75     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9701_5 ( .OUT(na9701_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2851_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9702_5 ( .OUT(na9702_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2857_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9703_5 ( .OUT(na9703_2), .IN1(1'b0), .IN2(na2894_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y105     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9704_5 ( .OUT(na9704_2), .IN1(1'b0), .IN2(na2895_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y49     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9705_5 ( .OUT(na9705_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2907_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y82     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9706_5 ( .OUT(na9706_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2908_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9707_5 ( .OUT(na9707_2), .IN1(1'b0), .IN2(na2910_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x130y80     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9708_5 ( .OUT(na9708_2), .IN1(1'b0), .IN2(na2911_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y84     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9709_5 ( .OUT(na9709_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2912_1), .IN8(1'b0) );
// C_////Bridge      x123y86     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9710_5 ( .OUT(na9710_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2913_1) );
// C_////Bridge      x127y89     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9711_5 ( .OUT(na9711_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2914_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y85     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9712_5 ( .OUT(na9712_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2915_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y104     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9713_5 ( .OUT(na9713_2), .IN1(1'b0), .IN2(na2919_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9714_5 ( .OUT(na9714_2), .IN1(1'b0), .IN2(na2935_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y94     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9715_5 ( .OUT(na9715_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2937_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y82     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9716_5 ( .OUT(na9716_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2943_1) );
// C_////Bridge      x127y87     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9717_5 ( .OUT(na9717_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2944_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9718_5 ( .OUT(na9718_2), .IN1(1'b0), .IN2(na2945_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9719_5 ( .OUT(na9719_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2953_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x127y75     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9720_5 ( .OUT(na9720_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2955_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y77     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9721_5 ( .OUT(na9721_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2957_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9722_5 ( .OUT(na9722_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2966_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y75     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9723_5 ( .OUT(na9723_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2967_1) );
// C_////Bridge      x90y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9724_5 ( .OUT(na9724_2), .IN1(1'b0), .IN2(na2971_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x130y48     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9725_5 ( .OUT(na9725_2), .IN1(1'b0), .IN2(na2972_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y38     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9726_5 ( .OUT(na9726_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2972_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9727_5 ( .OUT(na9727_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2974_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y89     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9728_5 ( .OUT(na9728_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2977_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9729_5 ( .OUT(na9729_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2979_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x120y47     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9730_5 ( .OUT(na9730_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2991_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y60     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9731_5 ( .OUT(na9731_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2995_1), .IN8(1'b0) );
// C_////Bridge      x99y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9732_5 ( .OUT(na9732_2), .IN1(na2996_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y78     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9733_5 ( .OUT(na9733_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3008_1) );
// C_////Bridge      x124y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9734_5 ( .OUT(na9734_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3010_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9735_5 ( .OUT(na9735_2), .IN1(1'b0), .IN2(na3011_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9736_5 ( .OUT(na9736_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3017_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x128y83     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9737_5 ( .OUT(na9737_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3017_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y46     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9738_5 ( .OUT(na9738_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3032_1) );
// C_////Bridge      x124y79     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9739_5 ( .OUT(na9739_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3066_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y95     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9740_5 ( .OUT(na9740_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3070_1) );
// C_////Bridge      x121y99     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9741_5 ( .OUT(na9741_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3071_1) );
// C_////Bridge      x115y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9742_5 ( .OUT(na9742_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3072_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9743_5 ( .OUT(na9743_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3072_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y97     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9744_5 ( .OUT(na9744_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3073_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9745_5 ( .OUT(na9745_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3073_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y94     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9746_5 ( .OUT(na9746_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3074_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y93     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9747_5 ( .OUT(na9747_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3075_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y87     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9748_5 ( .OUT(na9748_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3076_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x124y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9749_5 ( .OUT(na9749_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3076_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9750_5 ( .OUT(na9750_2), .IN1(1'b0), .IN2(na3107_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y84     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9751_5 ( .OUT(na9751_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3107_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x126y94     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9752_5 ( .OUT(na9752_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3110_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y91     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9753_5 ( .OUT(na9753_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3111_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y84     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9754_5 ( .OUT(na9754_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3116_1), .IN8(1'b0) );
// C_////Bridge      x90y99     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9755_5 ( .OUT(na9755_2), .IN1(na3118_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x122y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9756_5 ( .OUT(na9756_2), .IN1(na3121_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x125y93     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9757_5 ( .OUT(na9757_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3123_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9758_5 ( .OUT(na9758_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3124_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x118y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9759_5 ( .OUT(na9759_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3124_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y108     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9760_5 ( .OUT(na9760_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3126_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y89     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9761_5 ( .OUT(na9761_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3128_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y94     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9762_5 ( .OUT(na9762_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3128_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y91     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9763_5 ( .OUT(na9763_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3129_1) );
// C_////Bridge      x99y105     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9764_5 ( .OUT(na9764_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3130_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y80     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9765_5 ( .OUT(na9765_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3136_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y95     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9766_5 ( .OUT(na9766_2), .IN1(1'b0), .IN2(na3138_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y98     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9767_5 ( .OUT(na9767_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3141_1), .IN8(1'b0) );
// C_////Bridge      x98y93     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9768_5 ( .OUT(na9768_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3148_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y101     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9769_5 ( .OUT(na9769_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3151_1) );
// C_////Bridge      x109y93     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9770_5 ( .OUT(na9770_2), .IN1(1'b0), .IN2(na3152_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y101     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9771_5 ( .OUT(na9771_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3153_1) );
// C_////Bridge      x113y55     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9772_5 ( .OUT(na9772_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3154_1) );
// C_////Bridge      x119y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9773_5 ( .OUT(na9773_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3155_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9774_5 ( .OUT(na9774_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3155_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9775_5 ( .OUT(na9775_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3163_1) );
// C_////Bridge      x115y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9776_5 ( .OUT(na9776_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3164_1) );
// C_////Bridge      x98y102     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9777_5 ( .OUT(na9777_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3169_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y105     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9778_5 ( .OUT(na9778_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3170_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9779_5 ( .OUT(na9779_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3175_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x134y83     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9780_5 ( .OUT(na9780_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3175_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9781_5 ( .OUT(na9781_2), .IN1(1'b0), .IN2(na3178_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y64     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9782_5 ( .OUT(na9782_2), .IN1(na3180_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x113y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9783_5 ( .OUT(na9783_2), .IN1(na3180_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y97     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9784_5 ( .OUT(na9784_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3183_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9785_5 ( .OUT(na9785_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3183_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y59     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9786_5 ( .OUT(na9786_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3185_1) );
// C_////Bridge      x117y98     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9787_5 ( .OUT(na9787_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3189_1) );
// C_////Bridge      x96y96     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9788_5 ( .OUT(na9788_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3190_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y99     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9789_5 ( .OUT(na9789_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3200_1), .IN8(1'b0) );
// C_////Bridge      x118y102     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9790_5 ( .OUT(na9790_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3203_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y107     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9791_5 ( .OUT(na9791_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3205_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y106     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9792_5 ( .OUT(na9792_2), .IN1(na3208_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y83     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9793_5 ( .OUT(na9793_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3212_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9794_5 ( .OUT(na9794_2), .IN1(1'b0), .IN2(na3213_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y94     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9795_5 ( .OUT(na9795_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3216_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y65     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9796_5 ( .OUT(na9796_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3219_1), .IN8(1'b0) );
// C_////Bridge      x115y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9797_5 ( .OUT(na9797_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3219_2), .IN8(1'b0) );
// C_////Bridge      x122y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9798_5 ( .OUT(na9798_2), .IN1(1'b0), .IN2(na3222_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9799_5 ( .OUT(na9799_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3226_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y66     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9800_5 ( .OUT(na9800_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3226_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9801_5 ( .OUT(na9801_2), .IN1(na3256_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y62     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9802_5 ( .OUT(na9802_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3263_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y73     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9803_5 ( .OUT(na9803_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3264_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9804_5 ( .OUT(na9804_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3265_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9805_5 ( .OUT(na9805_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3266_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9806_5 ( .OUT(na9806_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3268_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9807_5 ( .OUT(na9807_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3269_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9808_5 ( .OUT(na9808_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3272_2) );
// C_////Bridge      x91y97     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9809_5 ( .OUT(na9809_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3276_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x114y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9810_5 ( .OUT(na9810_2), .IN1(na3290_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9811_5 ( .OUT(na9811_2), .IN1(na3290_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y92     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9812_5 ( .OUT(na9812_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3297_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9813_5 ( .OUT(na9813_2), .IN1(1'b0), .IN2(na3299_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9814_5 ( .OUT(na9814_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3301_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9815_5 ( .OUT(na9815_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3309_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9816_5 ( .OUT(na9816_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3309_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9817_5 ( .OUT(na9817_2), .IN1(na3313_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y104     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9818_5 ( .OUT(na9818_2), .IN1(na3313_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y82     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9819_5 ( .OUT(na9819_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3326_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y86     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9820_5 ( .OUT(na9820_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3329_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y72     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9821_5 ( .OUT(na9821_2), .IN1(1'b0), .IN2(na3330_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x116y70     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9822_5 ( .OUT(na9822_2), .IN1(1'b0), .IN2(na3345_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y117     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9823_5 ( .OUT(na9823_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3357_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y59     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9824_5 ( .OUT(na9824_2), .IN1(1'b0), .IN2(na3489_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y61     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9825_5 ( .OUT(na9825_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3491_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9826_5 ( .OUT(na9826_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3491_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y81     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9827_5 ( .OUT(na9827_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3562_1) );
// C_////Bridge      x91y92     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9828_5 ( .OUT(na9828_2), .IN1(na3588_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x121y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9829_5 ( .OUT(na9829_2), .IN1(na3594_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9830_5 ( .OUT(na9830_2), .IN1(na3594_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x117y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9831_5 ( .OUT(na9831_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3596_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y120     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9832_5 ( .OUT(na9832_2), .IN1(1'b0), .IN2(na3600_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y86     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9833_5 ( .OUT(na9833_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3610_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y52     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9834_5 ( .OUT(na9834_2), .IN1(na3621_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y61     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9835_5 ( .OUT(na9835_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3703_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9836_5 ( .OUT(na9836_2), .IN1(1'b0), .IN2(na3705_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y69     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9837_5 ( .OUT(na9837_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3707_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y70     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9838_5 ( .OUT(na9838_2), .IN1(1'b0), .IN2(na3709_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y68     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9839_5 ( .OUT(na9839_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3709_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y67     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9840_5 ( .OUT(na9840_2), .IN1(na3711_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y57     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9841_5 ( .OUT(na9841_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3711_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y64     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9842_5 ( .OUT(na9842_2), .IN1(1'b0), .IN2(na3712_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y62     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9843_5 ( .OUT(na9843_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3712_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9844_5 ( .OUT(na9844_2), .IN1(1'b0), .IN2(na3714_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9845_5 ( .OUT(na9845_2), .IN1(1'b0), .IN2(na3714_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y63     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9846_5 ( .OUT(na9846_2), .IN1(na3716_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y62     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9847_5 ( .OUT(na9847_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3718_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9848_5 ( .OUT(na9848_2), .IN1(na3720_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y59     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9849_5 ( .OUT(na9849_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3727_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y58     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9850_5 ( .OUT(na9850_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3727_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y62     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9851_5 ( .OUT(na9851_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3729_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y57     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9852_5 ( .OUT(na9852_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3731_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y68     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9853_5 ( .OUT(na9853_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3805_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y76     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9854_5 ( .OUT(na9854_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3941_1), .IN8(1'b0) );
// C_////Bridge      x78y83     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9855_5 ( .OUT(na9855_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3943_1) );
// C_////Bridge      x77y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9856_5 ( .OUT(na9856_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3954_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y88     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9857_5 ( .OUT(na9857_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3961_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9858_5 ( .OUT(na9858_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3963_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9859_5 ( .OUT(na9859_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3965_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x129y80     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9860_5 ( .OUT(na9860_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3975_1) );
// C_////Bridge      x131y78     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9861_5 ( .OUT(na9861_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3975_2) );
// C_////Bridge      x118y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9862_5 ( .OUT(na9862_2), .IN1(1'b0), .IN2(na4173_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y82     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9863_5 ( .OUT(na9863_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na4175_2), .IN8(1'b0) );
// C_////Bridge      x111y80     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9864_5 ( .OUT(na9864_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4894_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9865_5 ( .OUT(na9865_2), .IN1(na5229_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y62     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9866_5 ( .OUT(na9866_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5230_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y57     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9867_5 ( .OUT(na9867_2), .IN1(na5236_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9868_5 ( .OUT(na9868_2), .IN1(na5236_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9869_5 ( .OUT(na9869_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5237_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9870_5 ( .OUT(na9870_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5237_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9871_5 ( .OUT(na9871_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5238_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y79     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9872_5 ( .OUT(na9872_2), .IN1(na5239_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y55     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9873_5 ( .OUT(na9873_2), .IN1(na5240_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y69     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9874_5 ( .OUT(na9874_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5241_1), .IN8(1'b0) );
// C_////Bridge      x50y45     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9875_5 ( .OUT(na9875_2), .IN1(na5242_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9876_5 ( .OUT(na9876_2), .IN1(na5242_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y42     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9877_5 ( .OUT(na9877_2), .IN1(na5243_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y66     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9878_5 ( .OUT(na9878_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na5244_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9879_5 ( .OUT(na9879_2), .IN1(na5249_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y58     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9880_5 ( .OUT(na9880_2), .IN1(1'b0), .IN2(na5250_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y38     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9881_5 ( .OUT(na9881_2), .IN1(na5251_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y57     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9882_5 ( .OUT(na9882_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5252_1), .IN8(1'b0) );
// C_////Bridge      x50y39     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9883_5 ( .OUT(na9883_2), .IN1(na5253_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y59     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9884_5 ( .OUT(na9884_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5254_2), .IN8(1'b0) );
// C_////Bridge      x75y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9885_5 ( .OUT(na9885_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5255_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y71     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9886_5 ( .OUT(na9886_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5256_1), .IN8(1'b0) );
// C_////Bridge      x65y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9887_5 ( .OUT(na9887_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5257_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9888_5 ( .OUT(na9888_2), .IN1(1'b0), .IN2(na5258_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y37     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9889_5 ( .OUT(na9889_2), .IN1(na5259_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9890_5 ( .OUT(na9890_2), .IN1(na5261_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9891_5 ( .OUT(na9891_2), .IN1(1'b0), .IN2(na5266_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9892_5 ( .OUT(na9892_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5267_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9893_5 ( .OUT(na9893_2), .IN1(1'b0), .IN2(na5275_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y67     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9894_5 ( .OUT(na9894_2), .IN1(1'b0), .IN2(na5276_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9895_5 ( .OUT(na9895_2), .IN1(1'b0), .IN2(na5277_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9896_5 ( .OUT(na9896_2), .IN1(1'b0), .IN2(na5278_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y77     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9897_5 ( .OUT(na9897_2), .IN1(1'b0), .IN2(na5279_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9898_5 ( .OUT(na9898_2), .IN1(1'b0), .IN2(na5281_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y72     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9899_5 ( .OUT(na9899_2), .IN1(1'b0), .IN2(na5282_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9900_5 ( .OUT(na9900_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na5283_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9901_5 ( .OUT(na9901_2), .IN1(1'b0), .IN2(na5284_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9902_5 ( .OUT(na9902_2), .IN1(1'b0), .IN2(na5290_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9903_5 ( .OUT(na9903_2), .IN1(1'b0), .IN2(na5291_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y97     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9904_5 ( .OUT(na9904_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5435_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y68     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9905_5 ( .OUT(na9905_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5691_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9906_5 ( .OUT(na9906_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5691_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y57     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9907_5 ( .OUT(na9907_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5692_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9908_5 ( .OUT(na9908_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5705_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y53     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9909_5 ( .OUT(na9909_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na5705_2) );
// C_////Bridge      x75y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9910_5 ( .OUT(na9910_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5842_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9911_5 ( .OUT(na9911_2), .IN1(1'b0), .IN2(na5953_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y82     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9912_5 ( .OUT(na9912_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na5953_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y78     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9913_5 ( .OUT(na9913_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5955_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9914_5 ( .OUT(na9914_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5958_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9915_5 ( .OUT(na9915_2), .IN1(1'b0), .IN2(na5959_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y90     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9916_5 ( .OUT(na9916_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5961_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9917_5 ( .OUT(na9917_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5962_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9918_5 ( .OUT(na9918_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5962_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y90     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9919_5 ( .OUT(na9919_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5963_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y55     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9920_5 ( .OUT(na9920_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5964_1), .IN8(1'b0) );
// C_////Bridge      x55y53     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9921_5 ( .OUT(na9921_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5964_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y59     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9922_5 ( .OUT(na9922_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5965_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y61     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9923_5 ( .OUT(na9923_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5965_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9924_5 ( .OUT(na9924_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5967_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y50     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9925_5 ( .OUT(na9925_2), .IN1(na5967_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9926_5 ( .OUT(na9926_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5969_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y94     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9927_5 ( .OUT(na9927_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5969_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9928_5 ( .OUT(na9928_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5969_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y92     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9929_5 ( .OUT(na9929_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5969_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y91     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9930_5 ( .OUT(na9930_2), .IN1(na5971_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y56     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9931_5 ( .OUT(na9931_2), .IN1(na5971_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9932_5 ( .OUT(na9932_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na5971_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y48     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9933_5 ( .OUT(na9933_2), .IN1(na5972_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x136y115     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9934_5 ( .OUT(na9934_2), .IN1(na6055_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x123y111     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9935_5 ( .OUT(na9935_2), .IN1(1'b0), .IN2(na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9936_5 ( .OUT(na9936_2), .IN1(1'b0), .IN2(na6065_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9937_5 ( .OUT(na9937_2), .IN1(1'b0), .IN2(1'b0), .IN3(na6308_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9938_5 ( .OUT(na9938_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na6309_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y65     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9939_5 ( .OUT(na9939_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na6310_1) );
// C_////Bridge      x103y93     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9940_5 ( .OUT(na9940_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x119y60     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9941_5 ( .OUT(na9941_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9942_5 ( .OUT(na9942_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na6626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y93     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9943_5 ( .OUT(na9943_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na6661_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9944_5 ( .OUT(na9944_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na6673_1) );
// C_////Bridge      x105y62     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9945_5 ( .OUT(na9945_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na6673_2) );
// C_////Bridge      x93y70     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9946_5 ( .OUT(na9946_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na6675_2), .IN8(1'b0) );
// C_////Bridge      x99y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9947_5 ( .OUT(na9947_2), .IN1(1'b0), .IN2(1'b0), .IN3(na6684_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9948_5 ( .OUT(na9948_2), .IN1(1'b0), .IN2(1'b0), .IN3(na6684_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y90     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9949_5 ( .OUT(na9949_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na6727_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y48     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9950_5 ( .OUT(na9950_2), .IN1(1'b0), .IN2(1'b0), .IN3(na6947_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9951_5 ( .OUT(na9951_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7066_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9952_5 ( .OUT(na9952_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7112_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9953_5 ( .OUT(na9953_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7166_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y83     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9954_5 ( .OUT(na9954_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7210_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y64     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9955_5 ( .OUT(na9955_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7311_2), .IN8(1'b0) );
// C_////Bridge      x85y54     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9956_5 ( .OUT(na9956_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7411_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y54     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9957_5 ( .OUT(na9957_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7450_2), .IN8(1'b0) );
// C_////Bridge      x84y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9958_5 ( .OUT(na9958_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7495_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9959_5 ( .OUT(na9959_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7532_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y59     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9960_5 ( .OUT(na9960_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7567_2) );
// C_////Bridge      x57y59     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9961_5 ( .OUT(na9961_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7568_1) );
// C_////Bridge      x53y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9962_5 ( .OUT(na9962_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7570_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y61     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9963_5 ( .OUT(na9963_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7571_1), .IN8(1'b0) );
// C_////Bridge      x47y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9964_5 ( .OUT(na9964_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7572_2) );
// C_////Bridge      x49y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9965_5 ( .OUT(na9965_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7574_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y65     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9966_5 ( .OUT(na9966_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7575_2), .IN8(1'b0) );
// C_////Bridge      x53y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9967_5 ( .OUT(na9967_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7576_1), .IN8(1'b0) );
// C_////Bridge      x49y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9968_5 ( .OUT(na9968_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7578_2) );
// C_////Bridge      x49y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9969_5 ( .OUT(na9969_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7579_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y71     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9970_5 ( .OUT(na9970_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7580_2), .IN8(1'b0) );
// C_////Bridge      x47y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9971_5 ( .OUT(na9971_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7582_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9972_5 ( .OUT(na9972_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7583_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9973_5 ( .OUT(na9973_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7584_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9974_5 ( .OUT(na9974_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7586_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9975_5 ( .OUT(na9975_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7587_1), .IN8(1'b0) );
// C_////Bridge      x67y49     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9976_5 ( .OUT(na9976_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7588_2) );
// C_////Bridge      x73y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9977_5 ( .OUT(na9977_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7590_1) );
// C_////Bridge      x59y53     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9978_5 ( .OUT(na9978_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7591_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y53     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9979_5 ( .OUT(na9979_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7592_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y53     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9980_5 ( .OUT(na9980_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7801_2) );
// C_////Bridge      x80y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9981_5 ( .OUT(na9981_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7803_1) );
// C_////Bridge      x82y53     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9982_5 ( .OUT(na9982_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7813_2) );
// C_////Bridge      x80y49     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9983_5 ( .OUT(na9983_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7815_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y54     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9984_5 ( .OUT(na9984_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7827_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y56     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9985_5 ( .OUT(na9985_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7831_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9986_5 ( .OUT(na9986_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7835_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9987_5 ( .OUT(na9987_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7839_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y56     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9988_5 ( .OUT(na9988_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7843_2) );
// C_////Bridge      x83y62     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9989_5 ( .OUT(na9989_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7847_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9990_5 ( .OUT(na9990_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7851_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9991_5 ( .OUT(na9991_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7855_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y54     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9992_5 ( .OUT(na9992_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7859_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9993_5 ( .OUT(na9993_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7863_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9994_5 ( .OUT(na9994_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7867_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9995_5 ( .OUT(na9995_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7871_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y54     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9996_5 ( .OUT(na9996_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7875_2) );
// C_////Bridge      x53y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9997_5 ( .OUT(na9997_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7879_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9998_5 ( .OUT(na9998_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7883_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a9999_5 ( .OUT(na9999_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7887_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y50     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10000_5 ( .OUT(na10000_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7892_2) );
// C_////Bridge      x73y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10001_5 ( .OUT(na10001_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7894_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10002_5 ( .OUT(na10002_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7896_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10003_5 ( .OUT(na10003_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7898_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y39     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10004_5 ( .OUT(na10004_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7900_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y43     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10005_5 ( .OUT(na10005_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7902_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10006_5 ( .OUT(na10006_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7904_2), .IN8(1'b0) );
// C_////Bridge      x63y53     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10007_5 ( .OUT(na10007_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7906_1), .IN8(1'b0) );
// C_////Bridge      x59y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10008_5 ( .OUT(na10008_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7907_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10009_5 ( .OUT(na10009_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7908_1) );
// C_////Bridge      x61y53     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10010_5 ( .OUT(na10010_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7909_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10011_5 ( .OUT(na10011_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7911_1), .IN8(1'b0) );
// C_////Bridge      x65y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10012_5 ( .OUT(na10012_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7913_2) );
// C_////Bridge      x61y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10013_5 ( .OUT(na10013_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7914_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10014_5 ( .OUT(na10014_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na7915_2), .IN8(1'b0) );
// C_////Bridge      x63y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10015_5 ( .OUT(na10015_2), .IN1(1'b0), .IN2(1'b0), .IN3(na7916_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y45     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10016_5 ( .OUT(na10016_2), .IN1(na7966_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10017_5 ( .OUT(na10017_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8022_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10018_5 ( .OUT(na10018_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8023_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10019_5 ( .OUT(na10019_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8028_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y64     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10020_5 ( .OUT(na10020_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8029_1), .IN8(1'b0) );
// C_////Bridge      x82y50     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10021_5 ( .OUT(na10021_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8034_2), .IN8(1'b0) );
// C_////Bridge      x80y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10022_5 ( .OUT(na10022_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8035_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10023_5 ( .OUT(na10023_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8040_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10024_5 ( .OUT(na10024_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8041_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10025_5 ( .OUT(na10025_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8042_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10026_5 ( .OUT(na10026_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8043_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x115y75     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10027_5 ( .OUT(na10027_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8101_2), .IN8(1'b0) );
// C_////Bridge      x122y54     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10028_5 ( .OUT(na10028_2), .IN1(na8107_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10029_5 ( .OUT(na10029_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8164_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10030_5 ( .OUT(na10030_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8165_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10031_5 ( .OUT(na10031_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8170_2) );
// C_////Bridge      x78y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10032_5 ( .OUT(na10032_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8171_1) );
// C_////Bridge      x76y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10033_5 ( .OUT(na10033_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8179_2) );
// C_////Bridge      x82y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10034_5 ( .OUT(na10034_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8180_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10035_5 ( .OUT(na10035_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8183_1) );
// C_////Bridge      x86y61     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10036_5 ( .OUT(na10036_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8189_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y59     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10037_5 ( .OUT(na10037_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8191_1) );
// C_////Bridge      x82y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10038_5 ( .OUT(na10038_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8195_2) );
// C_////Bridge      x76y61     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10039_5 ( .OUT(na10039_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8196_1) );
// C_////Bridge      x86y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10040_5 ( .OUT(na10040_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8203_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10041_5 ( .OUT(na10041_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8206_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10042_5 ( .OUT(na10042_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8207_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10043_5 ( .OUT(na10043_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8210_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10044_5 ( .OUT(na10044_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8211_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10045_5 ( .OUT(na10045_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8214_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10046_5 ( .OUT(na10046_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8215_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10047_5 ( .OUT(na10047_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8218_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10048_5 ( .OUT(na10048_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8219_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y55     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10049_5 ( .OUT(na10049_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8285_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y38     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10050_5 ( .OUT(na10050_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8287_2), .IN8(1'b0) );
// C_////Bridge      x59y45     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10051_5 ( .OUT(na10051_2), .IN1(1'b0), .IN2(na8292_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y58     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10052_5 ( .OUT(na10052_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8302_2) );
// C_////Bridge      x82y77     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10053_5 ( .OUT(na10053_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8349_2) );
// C_////Bridge      x81y90     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10054_5 ( .OUT(na10054_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8373_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10055_5 ( .OUT(na10055_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8380_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y50     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10056_5 ( .OUT(na10056_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8381_1), .IN8(1'b0) );
// C_////Bridge      x134y107     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10057_5 ( .OUT(na10057_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na8394_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10058_5 ( .OUT(na10058_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8499_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10059_5 ( .OUT(na10059_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8500_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y68     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10060_5 ( .OUT(na10060_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8503_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y74     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10061_5 ( .OUT(na10061_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8504_1), .IN8(1'b0) );
// C_////Bridge      x50y72     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10062_5 ( .OUT(na10062_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8507_2), .IN8(1'b0) );
// C_////Bridge      x52y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10063_5 ( .OUT(na10063_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8508_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y52     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10064_5 ( .OUT(na10064_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8511_2), .IN8(1'b0) );
// C_////Bridge      x56y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10065_5 ( .OUT(na10065_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8512_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y75     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10066_5 ( .OUT(na10066_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8589_2) );
// C_////Bridge      x52y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10067_5 ( .OUT(na10067_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8590_1) );
// C_////Bridge      x52y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10068_5 ( .OUT(na10068_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8593_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10069_5 ( .OUT(na10069_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8594_1) );
// C_////Bridge      x54y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10070_5 ( .OUT(na10070_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8597_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10071_5 ( .OUT(na10071_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8598_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10072_5 ( .OUT(na10072_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8601_2) );
// C_////Bridge      x74y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10073_5 ( .OUT(na10073_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8602_1) );
// C_////Bridge      x59y42     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10074_5 ( .OUT(na10074_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8605_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y44     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10075_5 ( .OUT(na10075_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8606_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10076_5 ( .OUT(na10076_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8607_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10077_5 ( .OUT(na10077_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8608_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10078_5 ( .OUT(na10078_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8609_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y54     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10079_5 ( .OUT(na10079_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8610_1) );
// C_////Bridge      x57y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10080_5 ( .OUT(na10080_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8611_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y50     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10081_5 ( .OUT(na10081_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8612_1), .IN8(1'b0) );
// C_////Bridge      x65y50     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10082_5 ( .OUT(na10082_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8613_2) );
// C_////Bridge      x59y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10083_5 ( .OUT(na10083_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8614_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10084_5 ( .OUT(na10084_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8615_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10085_5 ( .OUT(na10085_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8616_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y60     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10086_5 ( .OUT(na10086_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8617_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y60     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10087_5 ( .OUT(na10087_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8618_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y60     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10088_5 ( .OUT(na10088_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8619_2), .IN8(1'b0) );
// C_////Bridge      x59y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10089_5 ( .OUT(na10089_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8620_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y76     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10090_5 ( .OUT(na10090_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8621_2) );
// C_////Bridge      x53y74     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10091_5 ( .OUT(na10091_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8622_1) );
// C_////Bridge      x47y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10092_5 ( .OUT(na10092_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8623_2), .IN8(1'b0) );
// C_////Bridge      x49y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10093_5 ( .OUT(na10093_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8624_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y72     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10094_5 ( .OUT(na10094_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8625_2) );
// C_////Bridge      x53y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10095_5 ( .OUT(na10095_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8626_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10096_5 ( .OUT(na10096_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8627_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10097_5 ( .OUT(na10097_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8628_1), .IN8(1'b0) );
// C_////Bridge      x66y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10098_5 ( .OUT(na10098_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8739_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10099_5 ( .OUT(na10099_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8740_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y39     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10100_5 ( .OUT(na10100_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8741_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y41     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10101_5 ( .OUT(na10101_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8742_1) );
// C_////Bridge      x58y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10102_5 ( .OUT(na10102_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8745_2) );
// C_////Bridge      x70y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10103_5 ( .OUT(na10103_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8746_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y49     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10104_5 ( .OUT(na10104_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8749_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y49     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10105_5 ( .OUT(na10105_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8750_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10106_5 ( .OUT(na10106_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8753_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y59     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10107_5 ( .OUT(na10107_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8754_1) );
// C_////Bridge      x79y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10108_5 ( .OUT(na10108_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8821_2) );
// C_////Bridge      x75y65     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10109_5 ( .OUT(na10109_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8822_1) );
// C_////Bridge      x79y65     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10110_5 ( .OUT(na10110_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8823_2), .IN8(1'b0) );
// C_////Bridge      x83y55     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10111_5 ( .OUT(na10111_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8824_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10112_5 ( .OUT(na10112_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8825_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10113_5 ( .OUT(na10113_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8826_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10114_5 ( .OUT(na10114_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8827_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y47     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10115_5 ( .OUT(na10115_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8828_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10116_5 ( .OUT(na10116_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8829_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y49     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10117_5 ( .OUT(na10117_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8830_1) );
// C_////Bridge      x79y55     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10118_5 ( .OUT(na10118_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8831_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y59     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10119_5 ( .OUT(na10119_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8832_1), .IN8(1'b0) );
// C_////Bridge      x54y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10120_5 ( .OUT(na10120_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8835_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10121_5 ( .OUT(na10121_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8836_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10122_5 ( .OUT(na10122_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8839_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10123_5 ( .OUT(na10123_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8840_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10124_5 ( .OUT(na10124_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8909_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y59     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10125_5 ( .OUT(na10125_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8910_1) );
// C_////Bridge      x87y55     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10126_5 ( .OUT(na10126_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8911_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y57     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10127_5 ( .OUT(na10127_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8912_1), .IN8(1'b0) );
// C_////Bridge      x81y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10128_5 ( .OUT(na10128_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8913_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10129_5 ( .OUT(na10129_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8914_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y55     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10130_5 ( .OUT(na10130_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8915_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10131_5 ( .OUT(na10131_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8916_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10132_5 ( .OUT(na10132_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8917_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10133_5 ( .OUT(na10133_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8918_1) );
// C_////Bridge      x75y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10134_5 ( .OUT(na10134_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8919_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y55     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10135_5 ( .OUT(na10135_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8920_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10136_5 ( .OUT(na10136_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8921_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10137_5 ( .OUT(na10137_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8922_1) );
// C_////Bridge      x79y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10138_5 ( .OUT(na10138_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8923_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10139_5 ( .OUT(na10139_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8924_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10140_5 ( .OUT(na10140_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8925_2) );
// C_////Bridge      x87y59     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10141_5 ( .OUT(na10141_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8926_1) );
// C_////Bridge      x87y65     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10142_5 ( .OUT(na10142_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8927_2), .IN8(1'b0) );
// C_////Bridge      x85y53     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10143_5 ( .OUT(na10143_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8928_1), .IN8(1'b0) );
// C_////Bridge      x75y64     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10144_5 ( .OUT(na10144_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8929_2) );
// C_////Bridge      x81y62     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10145_5 ( .OUT(na10145_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8930_1) );
// C_////Bridge      x75y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10146_5 ( .OUT(na10146_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8931_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10147_5 ( .OUT(na10147_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8932_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y62     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10148_5 ( .OUT(na10148_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8933_2) );
// C_////Bridge      x89y62     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10149_5 ( .OUT(na10149_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8934_1) );
// C_////Bridge      x89y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10150_5 ( .OUT(na10150_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8935_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10151_5 ( .OUT(na10151_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8936_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y66     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10152_5 ( .OUT(na10152_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8937_2) );
// C_////Bridge      x79y62     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10153_5 ( .OUT(na10153_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8938_1) );
// C_////Bridge      x73y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10154_5 ( .OUT(na10154_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8939_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10155_5 ( .OUT(na10155_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8940_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y52     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10156_5 ( .OUT(na10156_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8941_2) );
// C_////Bridge      x77y52     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10157_5 ( .OUT(na10157_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8942_1) );
// C_////Bridge      x81y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10158_5 ( .OUT(na10158_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8943_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y48     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10159_5 ( .OUT(na10159_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8944_1), .IN8(1'b0) );
// C_////Bridge      x81y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10160_5 ( .OUT(na10160_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na8945_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y50     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10161_5 ( .OUT(na10161_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na8946_1) );
// C_////Bridge      x85y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10162_5 ( .OUT(na10162_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8947_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y60     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10163_5 ( .OUT(na10163_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8948_1), .IN8(1'b0) );
// C_////Bridge      x97y85     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a10164_5 ( .OUT(na10164_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na9123_2), .IN8(1'b0) );
endmodule
